# 
# LEF OUT 
# User Name : m101jhwu 
# Date : Wed Nov 13 11:17:37 2013
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;

LAYER JX
  TYPE MASTERSLICE ;
END JX

LAYER RX
  TYPE MASTERSLICE ;
END RX

LAYER T3
  TYPE MASTERSLICE ;
END T3

LAYER NW
  TYPE MASTERSLICE ;
END NW

LAYER ALPHA
  TYPE MASTERSLICE ;
END ALPHA

LAYER PC
  TYPE MASTERSLICE ;
END PC

LAYER DG_BASE0
  TYPE MASTERSLICE ;
END DG_BASE0

LAYER CA
  TYPE MASTERSLICE ;
END CA

LAYER DV_BASE0
  TYPE MASTERSLICE ;
END DV_BASE0

LAYER OP
  TYPE MASTERSLICE ;
END OP

LAYER TAP
  TYPE MASTERSLICE ;
END TAP

LAYER OUTLINE_BASE0
  TYPE MASTERSLICE ;
END OUTLINE_BASE0

LAYER TEXT
  TYPE MASTERSLICE ;
END TEXT

LAYER W0_BASE0
  TYPE MASTERSLICE ;
END W0_BASE0

LAYER B1_BASE0
  TYPE MASTERSLICE ;
END B1_BASE0

LAYER W1_BASE0
  TYPE MASTERSLICE ;
END W1_BASE0

LAYER B2_BASE0
  TYPE MASTERSLICE ;
END B2_BASE0

LAYER W2_BASE0
  TYPE MASTERSLICE ;
END W2_BASE0

LAYER B3_BASE0
  TYPE MASTERSLICE ;
END B3_BASE0

LAYER W3_BASE0
  TYPE MASTERSLICE ;
END W3_BASE0

LAYER B4_BASE0
  TYPE MASTERSLICE ;
END B4_BASE0

LAYER WT_BASE0
  TYPE MASTERSLICE ;
END WT_BASE0

LAYER BA_BASE0
  TYPE MASTERSLICE ;
END BA_BASE0

LAYER WA_BASE0
  TYPE MASTERSLICE ;
END WA_BASE0

LAYER BB_BASE0
  TYPE MASTERSLICE ;
END BB_BASE0

LAYER WB_BASE0
  TYPE MASTERSLICE ;
END WB_BASE0

LAYER BD_BASE0
  TYPE MASTERSLICE ;
END BD_BASE0

LAYER WD_BASE0
  TYPE MASTERSLICE ;
END WD_BASE0

LAYER BE_BASE0
  TYPE MASTERSLICE ;
END BE_BASE0

LAYER YT_BASE0
  TYPE MASTERSLICE ;
END YT_BASE0

LAYER YA_BASE0
  TYPE MASTERSLICE ;
END YA_BASE0

LAYER EB_BASE0
  TYPE MASTERSLICE ;
END EB_BASE0

LAYER N3
  TYPE MASTERSLICE ;
END N3

LAYER BG
  TYPE MASTERSLICE ;
END BG

LAYER WE
  TYPE MASTERSLICE ;
END WE

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.09 ;
  OFFSET 0.1 ;
  AREA 0.042 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      0.38   0.42   1.5    4.5    
      WIDTH 0           0.09   0.11   0.16   0.5    1.5    
      WIDTH 0.2         0.11   0.11   0.16   0.5    1.5    
      WIDTH 0.42        0.16   0.16   0.16   0.5    1.5    
      WIDTH 1.5         0.5    0.5    0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    1.5    1.5    ;
  MAXWIDTH 12 ;
  MINWIDTH 0.09 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.122 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 25 25 ;
  DENSITYCHECKSTEP 12.5 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.13 ;
  SPACING 0 ADJACENTCUTS 3 WITHIN 0.14 ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      0.38   0.42   1.5    4.5    
      WIDTH 0           0.1    0.12   0.16   0.5    1.5    
      WIDTH 0.2         0.12   0.12   0.16   0.5    1.5    
      WIDTH 0.42        0.16   0.16   0.16   0.5    1.5    
      WIDTH 1.5         0.5    0.5    0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    1.5    1.5    ;
  MAXWIDTH 12 ;
  MINWIDTH 0.1 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.124 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.13 ;
  SPACING 0 ADJACENTCUTS 3 WITHIN 0.14 ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      0.38   0.42   1.5    4.5    
      WIDTH 0           0.1    0.12   0.16   0.5    1.5    
      WIDTH 0.2         0.12   0.12   0.16   0.5    1.5    
      WIDTH 0.42        0.16   0.16   0.16   0.5    1.5    
      WIDTH 1.5         0.5    0.5    0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    1.5    1.5    ;
  MAXWIDTH 12 ;
  MINWIDTH 0.1 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.124 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M3

LAYER V3
  TYPE CUT ;
  SPACING 0.13 ;
  SPACING 0 ADJACENTCUTS 3 WITHIN 0.14 ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      0.38   0.42   1.5    4.5    
      WIDTH 0           0.1    0.12   0.16   0.5    1.5    
      WIDTH 0.2         0.12   0.12   0.16   0.5    1.5    
      WIDTH 0.42        0.16   0.16   0.16   0.5    1.5    
      WIDTH 1.5         0.5    0.5    0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    1.5    1.5    ;
  MAXWIDTH 12 ;
  MINWIDTH 0.1 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.124 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M4

LAYER V4
  TYPE CUT ;
  SPACING 0.13 ;
  SPACING 0 ADJACENTCUTS 3 WITHIN 0.14 ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      0.38   0.42   1.5    4.5    
      WIDTH 0           0.1    0.12   0.16   0.5    1.5    
      WIDTH 0.2         0.12   0.12   0.16   0.5    1.5    
      WIDTH 0.42        0.16   0.16   0.16   0.5    1.5    
      WIDTH 1.5         0.5    0.5    0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    1.5    1.5    ;
  MAXWIDTH 12 ;
  MINWIDTH 0.1 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.124 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M5

LAYER V5
  TYPE CUT ;
  SPACING 0.13 ;
  SPACING 0 ADJACENTCUTS 3 WITHIN 0.14 ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      0.38   0.42   1.5    4.5    
      WIDTH 0           0.1    0.12   0.16   0.5    1.5    
      WIDTH 0.2         0.12   0.12   0.16   0.5    1.5    
      WIDTH 0.42        0.16   0.16   0.16   0.5    1.5    
      WIDTH 1.5         0.5    0.5    0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    1.5    1.5    ;
  MAXWIDTH 12 ;
  MINWIDTH 0.1 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.124 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M6

LAYER NT
  TYPE CUT ;
  SPACING 0.44 ;
  SPACING 0 ADJACENTCUTS 3 WITHIN 0.56 ;
END NT

LAYER EA
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.8 ;
  WIDTH 0.4 ;
  OFFSET 0.1 ;
  AREA 0.565 ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0      1.5    4.5    
      WIDTH 0           0.4    0.5    1.5    
      WIDTH 1.5         0.5    0.5    1.5    
      WIDTH 4.5         1.5    1.5    1.5    ;
  MINIMUMCUT 2 WIDTH 1.804 ;
  MAXWIDTH 12.25 ;
  MINWIDTH 0.4 ;
  MINENCLOSEDAREA 0.565 ;
  RESISTANCE RPERSQ 0.0279 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END EA

LAYER VV
  TYPE CUT ;
  SPACING 2 ;
END VV

LAYER LB
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 6 ;
  WIDTH 3 ;
  OFFSET 0.1 ;
  SPACING 2 ;
  MINIMUMCUT 2 WIDTH 1.804 ;
  MINWIDTH 3 ;
  RESISTANCE RPERSQ 0.0275 ;
  CAPMULTIPLIER 1 ;
END LB

LAYER OverlapCheck
  TYPE OVERLAP ;
END OverlapCheck

VIA V1_0_HH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_0_HH_F0

VIA V1_0_HH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_0_HH_F1

VIA V1_0_HV_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_0_HV_F0

VIA V1_0_HV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_0_HV_F1

VIA V1_0_VH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_0_VH_F0

VIA V1_0_VH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_0_VH_F1

VIA V1_0_VV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_0_VV_F0

VIA V1_0_VV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_0_VV_F1

VIA V1_1_HH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_1_HH_F0

VIA V1_1_HH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_1_HH_F1

VIA V1_1_HV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_1_HV_F0

VIA V1_1_HV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_1_HV_F1

VIA V1_1_VH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_1_VH_F0

VIA V1_1_VH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_1_VH_F1

VIA V1_1_VV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_1_VV_F0

VIA V1_1_VV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_1_VV_F1

VIA V1_2_XH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_2_XH_F0

VIA V1_2_XH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V1_2_XH_F1

VIA V1_2_XV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_2_XV_F0

VIA V1_2_XV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V1_2_XV_F1

VIA V1_3_HH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_3_HH_F0

VIA V1_3_HH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_3_HH_F1

VIA V1_3_HV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_3_HV_F0

VIA V1_3_HV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_3_HV_F1

VIA V1_3_VH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_3_VH_F0

VIA V1_3_VH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_3_VH_F1

VIA V1_3_VV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_3_VV_F0

VIA V1_3_VV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_3_VV_F1

VIA V1_4_HH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_4_HH_F0

VIA V1_4_HH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_4_HH_F1

VIA V1_4_HV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_4_HV_F0

VIA V1_4_HV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_4_HV_F1

VIA V1_4_VH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_4_VH_F0

VIA V1_4_VH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_4_VH_F1

VIA V1_4_VV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_4_VV_F0

VIA V1_4_VV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_4_VV_F1

VIA V1_5_XH_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_5_XH_F0

VIA V1_5_XH_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V1_5_XH_F1

VIA V1_5_XV_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_5_XV_F0

VIA V1_5_XV_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V1_5_XV_F1

VIA V1_6_HX_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_6_HX_F0

VIA V1_6_HX_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_6_HX_F1

VIA V1_6_VX_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_6_VX_F0

VIA V1_6_VX_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_6_VX_F1

VIA V1_7_HX_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_7_HX_F0

VIA V1_7_HX_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_7_HX_F1

VIA V1_7_VX_F0
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_7_VX_F0

VIA V1_7_VX_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_7_VX_F1

VIA V1_8_XX_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_8_XX_F0

VIA V1_8_XX_F1
  RESISTANCE 7 ;
  LAYER M1 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V1_8_XX_F1

VIA V2_0_HH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_0_HH_F0

VIA V2_0_HH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_0_HH_F1

VIA V2_0_HV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_0_HV_F0

VIA V2_0_HV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_0_HV_F1

VIA V2_0_VH_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_0_VH_F0

VIA V2_0_VH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_0_VH_F1

VIA V2_0_VV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_0_VV_F0

VIA V2_0_VV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_0_VV_F1

VIA V2_1_HH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_1_HH_F0

VIA V2_1_HH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_1_HH_F1

VIA V2_1_HV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_1_HV_F0

VIA V2_1_HV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_1_HV_F1

VIA V2_1_VH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_1_VH_F0

VIA V2_1_VH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_1_VH_F1

VIA V2_1_VV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_1_VV_F0

VIA V2_1_VV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_1_VV_F1

VIA V2_2_XH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_2_XH_F0

VIA V2_2_XH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V2_2_XH_F1

VIA V2_2_XV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_2_XV_F0

VIA V2_2_XV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V2_2_XV_F1

VIA V2_3_HH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_3_HH_F0

VIA V2_3_HH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_3_HH_F1

VIA V2_3_HV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_3_HV_F0

VIA V2_3_HV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_3_HV_F1

VIA V2_3_VH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_3_VH_F0

VIA V2_3_VH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_3_VH_F1

VIA V2_3_VV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_3_VV_F0

VIA V2_3_VV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_3_VV_F1

VIA V2_4_HH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_4_HH_F0

VIA V2_4_HH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_4_HH_F1

VIA V2_4_HV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_4_HV_F0

VIA V2_4_HV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_4_HV_F1

VIA V2_4_VH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_4_VH_F0

VIA V2_4_VH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_4_VH_F1

VIA V2_4_VV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_4_VV_F0

VIA V2_4_VV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_4_VV_F1

VIA V2_5_XH_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_5_XH_F0

VIA V2_5_XH_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V2_5_XH_F1

VIA V2_5_XV_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_5_XV_F0

VIA V2_5_XV_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V2_5_XV_F1

VIA V2_6_HX_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_6_HX_F0

VIA V2_6_HX_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_6_HX_F1

VIA V2_6_VX_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_6_VX_F0

VIA V2_6_VX_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_6_VX_F1

VIA V2_7_HX_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_7_HX_F0

VIA V2_7_HX_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_7_HX_F1

VIA V2_7_VX_F0
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_7_VX_F0

VIA V2_7_VX_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_7_VX_F1

VIA V2_8_XX_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_8_XX_F0

VIA V2_8_XX_F1
  RESISTANCE 7 ;
  LAYER M2 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V2_8_XX_F1

VIA V3_0_HV_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_0_HV_F0

VIA V3_0_HV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_0_HV_F1

VIA V3_0_VV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_0_VV_F0

VIA V3_0_VV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_0_VV_F1

VIA V3_1_HV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_1_HV_F0

VIA V3_1_HV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_1_HV_F1

VIA V3_1_VV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_1_VV_F0

VIA V3_1_VV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_1_VV_F1

VIA V3_2_XV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_2_XV_F0

VIA V3_2_XV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V3_2_XV_F1

VIA V3_3_HV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_3_HV_F0

VIA V3_3_HV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_3_HV_F1

VIA V3_3_VV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_3_VV_F0

VIA V3_3_VV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_3_VV_F1

VIA V3_4_HV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_4_HV_F0

VIA V3_4_HV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_4_HV_F1

VIA V3_4_VV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_4_VV_F0

VIA V3_4_VV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_4_VV_F1

VIA V3_5_XV_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_5_XV_F0

VIA V3_5_XV_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V3_5_XV_F1

VIA V3_6_HX_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_6_HX_F0

VIA V3_6_HX_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_6_HX_F1

VIA V3_6_VX_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_6_VX_F0

VIA V3_6_VX_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_6_VX_F1

VIA V3_7_HX_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_7_HX_F0

VIA V3_7_HX_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_7_HX_F1

VIA V3_7_VX_F0
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_7_VX_F0

VIA V3_7_VX_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_7_VX_F1

VIA V3_8_XX_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_8_XX_F0

VIA V3_8_XX_F1
  RESISTANCE 7 ;
  LAYER M3 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V3_8_XX_F1

VIA V4_0_VH_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V4_0_VH_F0

VIA V4_0_VH_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V4_0_VH_F1

VIA V4_1_VH_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V4_1_VH_F0

VIA V4_1_VH_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V4_1_VH_F1

VIA V4_2_XH_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V4_2_XH_F0

VIA V4_2_XH_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
END V4_2_XH_F1

VIA V4_3_VH_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V4_3_VH_F0

VIA V4_3_VH_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V4_3_VH_F1

VIA V4_4_VH_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V4_4_VH_F0

VIA V4_4_VH_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V4_4_VH_F1

VIA V4_5_XH_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V4_5_XH_F0

VIA V4_5_XH_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
END V4_5_XH_F1

VIA V4_6_VX_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V4_6_VX_F0

VIA V4_6_VX_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V4_6_VX_F1

VIA V4_7_VX_F0
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V4_7_VX_F0

VIA V4_7_VX_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V4_7_VX_F1

VIA V4_8_XX_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V4_8_XX_F0

VIA V4_8_XX_F1
  RESISTANCE 7 ;
  LAYER M4 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V4_8_XX_F1

VIA V5_0_HV_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V5_0_HV_F0

VIA V5_0_HV_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V5_0_HV_F1

VIA V5_1_HV_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V5_1_HV_F0

VIA V5_1_HV_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V5_1_HV_F1

VIA V5_2_XV_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V5_2_XV_F0

VIA V5_2_XV_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0500 -0.0900 0.0500 0.0900 ;
END V5_2_XV_F1

VIA V5_3_HV_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V5_3_HV_F0

VIA V5_3_HV_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V5_3_HV_F1

VIA V5_4_HV_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V5_4_HV_F0

VIA V5_4_HV_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V5_4_HV_F1

VIA V5_5_XV_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V5_5_XV_F0

VIA V5_5_XV_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0600 -0.0800 0.0600 0.0800 ;
END V5_5_XV_F1

VIA V5_6_HX_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V5_6_HX_F0

VIA V5_6_HX_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0900 -0.0500 0.0900 0.0500 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V5_6_HX_F1

VIA V5_7_HX_F0
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V5_7_HX_F0

VIA V5_7_HX_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0800 -0.0600 0.0800 0.0600 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V5_7_HX_F1

VIA V5_8_XX_F0
  DEFAULT 
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V5_8_XX_F0

VIA V5_8_XX_F1
  RESISTANCE 7 ;
  LAYER M5 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0700 -0.0700 0.0700 0.0700 ;
END V5_8_XX_F1

VIA NT_0_VH
  DEFAULT 
  RESISTANCE 1 ;
  LAYER M6 ;
    RECT -0.2000 -0.2600 0.2000 0.2600 ;
  LAYER NT ;
    RECT -0.1800 -0.1800 0.1800 0.1800 ;
  LAYER EA ;
    RECT -0.2600 -0.2000 0.2600 0.2000 ;
END NT_0_VH

VIA VV_0_HV
  DEFAULT 
  RESISTANCE 0.1 ;
  LAYER EA ;
    RECT -2.2500 -2.2500 2.2500 2.2500 ;
  LAYER VV ;
    RECT -1.5000 -1.5000 1.5000 1.5000 ;
  LAYER LB ;
    RECT -2.5000 -2.5000 2.5000 2.5000 ;
END VV_0_HV

VIARULE V1_0_HH_F0 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.04 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_HH_F0

VIARULE V1_0_HH_F1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.04 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_HH_F1

VIARULE V1_0_HV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_HV_F0

VIARULE V1_0_HV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_HV_F1

VIARULE V1_0_VH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_VH_F0

VIARULE V1_0_VH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_VH_F1

VIARULE V1_0_VV_F0 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_VV_F0

VIARULE V1_0_VV_F1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_0_VV_F1

VIARULE V1_1_HH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_HH_F0

VIARULE V1_1_HH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_HH_F1

VIARULE V1_1_HV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_HV_F0

VIARULE V1_1_HV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_HV_F1

VIARULE V1_1_VH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_VH_F0

VIARULE V1_1_VH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_VH_F1

VIARULE V1_1_VV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_VV_F0

VIARULE V1_1_VV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_1_VV_F1

VIARULE V1_2_XH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_2_XH_F0

VIARULE V1_2_XH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_2_XH_F1

VIARULE V1_2_XV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_2_XV_F0

VIARULE V1_2_XV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_2_XV_F1

VIARULE V1_3_HH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_HH_F0

VIARULE V1_3_HH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_HH_F1

VIARULE V1_3_HV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_HV_F0

VIARULE V1_3_HV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_HV_F1

VIARULE V1_3_VH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_VH_F0

VIARULE V1_3_VH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_VH_F1

VIARULE V1_3_VV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_VV_F0

VIARULE V1_3_VV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_3_VV_F1

VIARULE V1_4_HH_F0 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_HH_F0

VIARULE V1_4_HH_F1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_HH_F1

VIARULE V1_4_HV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_HV_F0

VIARULE V1_4_HV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_HV_F1

VIARULE V1_4_VH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_VH_F0

VIARULE V1_4_VH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_VH_F1

VIARULE V1_4_VV_F0 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_VV_F0

VIARULE V1_4_VV_F1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_4_VV_F1

VIARULE V1_5_XH_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_5_XH_F0

VIARULE V1_5_XH_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_5_XH_F1

VIARULE V1_5_XV_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_5_XV_F0

VIARULE V1_5_XV_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_5_XV_F1

VIARULE V1_6_HX_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_6_HX_F0

VIARULE V1_6_HX_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.04 0 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_6_HX_F1

VIARULE V1_6_VX_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_6_VX_F0

VIARULE V1_6_VX_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_6_VX_F1

VIARULE V1_7_HX_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_7_HX_F0

VIARULE V1_7_HX_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_7_HX_F1

VIARULE V1_7_VX_F0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_7_VX_F0

VIARULE V1_7_VX_F1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_7_VX_F1

VIARULE V1_8_XX_F0 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_8_XX_F0

VIARULE V1_8_XX_F1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER V1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V1_8_XX_F1

VIARULE V2_0_HH_F0 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_HH_F0

VIARULE V2_0_HH_F1 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_HH_F1

VIARULE V2_0_HV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_HV_F0

VIARULE V2_0_HV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_HV_F1

VIARULE V2_0_VH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_VH_F0

VIARULE V2_0_VH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_VH_F1

VIARULE V2_0_VV_F0 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.04 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_VV_F0

VIARULE V2_0_VV_F1 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.04 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_0_VV_F1

VIARULE V2_1_HH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_HH_F0

VIARULE V2_1_HH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_HH_F1

VIARULE V2_1_HV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_HV_F0

VIARULE V2_1_HV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_HV_F1

VIARULE V2_1_VH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_VH_F0

VIARULE V2_1_VH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_VH_F1

VIARULE V2_1_VV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_VV_F0

VIARULE V2_1_VV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_1_VV_F1

VIARULE V2_2_XH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_2_XH_F0

VIARULE V2_2_XH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_2_XH_F1

VIARULE V2_2_XV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_2_XV_F0

VIARULE V2_2_XV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_2_XV_F1

VIARULE V2_3_HH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_HH_F0

VIARULE V2_3_HH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_HH_F1

VIARULE V2_3_HV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_HV_F0

VIARULE V2_3_HV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_HV_F1

VIARULE V2_3_VH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_VH_F0

VIARULE V2_3_VH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_VH_F1

VIARULE V2_3_VV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_VV_F0

VIARULE V2_3_VV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_3_VV_F1

VIARULE V2_4_HH_F0 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_HH_F0

VIARULE V2_4_HH_F1 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.01 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_HH_F1

VIARULE V2_4_HV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_HV_F0

VIARULE V2_4_HV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_HV_F1

VIARULE V2_4_VH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_VH_F0

VIARULE V2_4_VH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_VH_F1

VIARULE V2_4_VV_F0 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_VV_F0

VIARULE V2_4_VV_F1 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_4_VV_F1

VIARULE V2_5_XH_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_5_XH_F0

VIARULE V2_5_XH_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_5_XH_F1

VIARULE V2_5_XV_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_5_XV_F0

VIARULE V2_5_XV_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_5_XV_F1

VIARULE V2_6_HX_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_6_HX_F0

VIARULE V2_6_HX_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.04 0 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_6_HX_F1

VIARULE V2_6_VX_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_6_VX_F0

VIARULE V2_6_VX_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_6_VX_F1

VIARULE V2_7_HX_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_7_HX_F0

VIARULE V2_7_HX_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_7_HX_F1

VIARULE V2_7_VX_F0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_7_VX_F0

VIARULE V2_7_VX_F1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_7_VX_F1

VIARULE V2_8_XX_F0 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_8_XX_F0

VIARULE V2_8_XX_F1 GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER V2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V2_8_XX_F1

VIARULE V3_0_HV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_0_HV_F0

VIARULE V3_0_HV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_0_HV_F1

VIARULE V3_0_VV_F0 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_0_VV_F0

VIARULE V3_0_VV_F1 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_0_VV_F1

VIARULE V3_1_HV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_1_HV_F0

VIARULE V3_1_HV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_1_HV_F1

VIARULE V3_1_VV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_1_VV_F0

VIARULE V3_1_VV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_1_VV_F1

VIARULE V3_2_XV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_2_XV_F0

VIARULE V3_2_XV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_2_XV_F1

VIARULE V3_3_HV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_3_HV_F0

VIARULE V3_3_HV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_3_HV_F1

VIARULE V3_3_VV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_3_VV_F0

VIARULE V3_3_VV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_3_VV_F1

VIARULE V3_4_HV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_4_HV_F0

VIARULE V3_4_HV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_4_HV_F1

VIARULE V3_4_VV_F0 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_4_VV_F0

VIARULE V3_4_VV_F1 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.01 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_4_VV_F1

VIARULE V3_5_XV_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_5_XV_F0

VIARULE V3_5_XV_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_5_XV_F1

VIARULE V3_6_HX_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_6_HX_F0

VIARULE V3_6_HX_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.04 0 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_6_HX_F1

VIARULE V3_6_VX_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_6_VX_F0

VIARULE V3_6_VX_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.04 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_6_VX_F1

VIARULE V3_7_HX_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_7_HX_F0

VIARULE V3_7_HX_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_7_HX_F1

VIARULE V3_7_VX_F0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_7_VX_F0

VIARULE V3_7_VX_F1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_7_VX_F1

VIARULE V3_8_XX_F0 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_8_XX_F0

VIARULE V3_8_XX_F1 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER V3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V3_8_XX_F1

VIARULE V4_0_VH_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_0_VH_F0

VIARULE V4_0_VH_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_0_VH_F1

VIARULE V4_1_VH_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_1_VH_F0

VIARULE V4_1_VH_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_1_VH_F1

VIARULE V4_2_XH_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_2_XH_F0

VIARULE V4_2_XH_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_2_XH_F1

VIARULE V4_3_VH_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_3_VH_F0

VIARULE V4_3_VH_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_3_VH_F1

VIARULE V4_4_VH_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_4_VH_F0

VIARULE V4_4_VH_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_4_VH_F1

VIARULE V4_5_XH_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_5_XH_F0

VIARULE V4_5_XH_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_5_XH_F1

VIARULE V4_6_VX_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_6_VX_F0

VIARULE V4_6_VX_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_6_VX_F1

VIARULE V4_7_VX_F0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_7_VX_F0

VIARULE V4_7_VX_F1 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_7_VX_F1

VIARULE V4_8_XX_F0 GENERATE
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_8_XX_F0

VIARULE V4_8_XX_F1 GENERATE
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER V4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V4_8_XX_F1

VIARULE V5_0_HV_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER M6 ;
    ENCLOSURE 0 0.04 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_0_HV_F0

VIARULE V5_0_HV_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER M6 ;
    ENCLOSURE 0 0.04 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_0_HV_F1

VIARULE V5_1_HV_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M6 ;
    ENCLOSURE 0 0.04 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_1_HV_F0

VIARULE V5_1_HV_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M6 ;
    ENCLOSURE 0 0.04 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_1_HV_F1

VIARULE V5_2_XV_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M6 ;
    ENCLOSURE 0 0.04 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_2_XV_F0

VIARULE V5_2_XV_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M6 ;
    ENCLOSURE 0 0.04 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_2_XV_F1

VIARULE V5_3_HV_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER M6 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_3_HV_F0

VIARULE V5_3_HV_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER M6 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_3_HV_F1

VIARULE V5_4_HV_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M6 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_4_HV_F0

VIARULE V5_4_HV_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M6 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_4_HV_F1

VIARULE V5_5_XV_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M6 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_5_XV_F0

VIARULE V5_5_XV_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER M6 ;
    ENCLOSURE 0.01 0.03 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_5_XV_F1

VIARULE V5_6_HX_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER M6 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_6_HX_F0

VIARULE V5_6_HX_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.04 0 ;
  LAYER M6 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_6_HX_F1

VIARULE V5_7_HX_F0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M6 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_7_HX_F0

VIARULE V5_7_HX_F1 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.01 ;
  LAYER M6 ;
    ENCLOSURE 0.02 0.02 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_7_HX_F1

VIARULE V5_8_XX_F0 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_8_XX_F0

VIARULE V5_8_XX_F1 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.02 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.02 ;
  LAYER V5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.23 BY 0.23 ;
    RESISTANCE 7 ;
END V5_8_XX_F1

VIARULE NT_0_VH GENERATE
  LAYER M6 ;
    ENCLOSURE 0.02 0.08 ;
  LAYER EA ;
    ENCLOSURE 0.08 0.02 ;
  LAYER NT ;
    RECT -0.1800 -0.1800 0.1800 0.1800 ;
    SPACING 0.8 BY 0.8 ;
    RESISTANCE 1 ;
END NT_0_VH

VIARULE VV_0_HV GENERATE
  LAYER EA ;
    ENCLOSURE 0.75 0.75 ;
  LAYER LB ;
    ENCLOSURE 1 1 ;
  LAYER VV ;
    RECT -1.5000 -1.5000 1.5000 1.5000 ;
    SPACING 5 BY 5 ;
    RESISTANCE 0.1 ;
END VV_0_HV

SPACING
  SAMENET V1 V1 0.1 ;
  SAMENET V2 V2 0.1 ;
  SAMENET V3 V3 0.1 ;
  SAMENET V4 V4 0.1 ;
  SAMENET V5 V5 0.1 ;
  SAMENET NT NT 0.34 ;
  SAMENET V2 V1 0 STACK ;
  SAMENET V3 V2 0 STACK ;
  SAMENET V4 V3 0 STACK ;
  SAMENET V5 V4 0 STACK ;
  SAMENET NT V5 0 STACK ;
END SPACING

SITE unit
  CLASS CORE ;
  SYMMETRY X Y ;
  SIZE 0.2 BY 2.4 ;
END unit

MACRO XOR3_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6150 ;
        RECT 3.2300 0.3200 3.4500 0.4050 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.7500 1.5500 ;
        RECT 0.6500 1.5500 0.7500 1.8200 ;
        RECT 0.2500 1.1400 0.3500 1.4500 ;
        RECT 0.6500 1.8200 1.5100 1.9200 ;
        RECT 0.2500 1.0400 0.9600 1.1400 ;
        RECT 1.3400 1.9200 1.5100 1.9850 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6300 0.5750 3.7500 1.8100 ;
    END
    ANTENNADIFFAREA 0.187275 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0350 0.8600 2.1500 1.8200 ;
        RECT 2.0350 1.8200 3.0100 1.9200 ;
    END
    ANTENNAGATEAREA 0.0879 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.2500 1.0000 1.3500 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 3.3250 1.7900 3.4950 2.0800 ;
        RECT 0.3900 1.7100 0.5000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2600 1.3300 2.3500 1.7200 ;
      RECT 2.2600 1.2400 2.5950 1.3300 ;
      RECT 2.5050 0.9700 2.5950 1.2400 ;
      RECT 2.2400 0.8800 2.5950 0.9700 ;
      RECT 2.2400 0.7500 2.3300 0.8800 ;
      RECT 2.0850 0.6600 2.3300 0.7500 ;
      RECT 0.8750 0.4800 2.5300 0.5700 ;
      RECT 2.4400 0.5700 2.5300 0.6800 ;
      RECT 2.4400 0.6800 2.8350 0.7700 ;
      RECT 2.7450 0.7700 2.8350 0.9150 ;
      RECT 2.7450 0.9150 3.1800 1.0050 ;
      RECT 2.7450 1.0050 2.8350 1.4300 ;
      RECT 2.5100 1.4300 2.8350 1.5200 ;
      RECT 2.5100 1.5200 2.6000 1.6550 ;
      RECT 1.1350 1.6400 1.8750 1.7300 ;
      RECT 1.7850 0.5700 1.8750 1.6400 ;
      RECT 3.0200 1.3950 3.3600 1.4850 ;
      RECT 3.2700 0.7700 3.3600 1.3950 ;
      RECT 2.9450 0.6800 3.3600 0.7700 ;
      RECT 2.7150 1.6100 3.5400 1.7000 ;
      RECT 3.4500 0.5900 3.5400 1.6100 ;
      RECT 2.6550 0.5000 3.5400 0.5900 ;
      RECT 0.0500 0.8400 1.1800 0.9300 ;
      RECT 1.0900 0.9300 1.1800 1.1450 ;
      RECT 0.0500 1.6600 0.2450 1.7500 ;
      RECT 0.0500 0.9300 0.1400 1.6600 ;
      RECT 0.0500 0.5050 0.1700 0.8400 ;
      RECT 0.9100 1.5450 1.0000 1.6800 ;
      RECT 0.9100 1.4550 1.4100 1.5450 ;
      RECT 1.3200 0.7500 1.4100 1.4550 ;
      RECT 0.6150 0.6600 1.4100 0.7500 ;
      RECT 1.5000 0.7500 1.5900 1.5300 ;
      RECT 1.5000 0.6600 1.6700 0.7500 ;
  END
END XOR3_X0P7M_A12TH

MACRO XOR3_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.8700 0.3500 1.3600 ;
        RECT 0.2450 0.7700 1.0400 0.8700 ;
        RECT 0.9400 0.8700 1.0400 1.0500 ;
        RECT 0.9400 1.0500 1.2600 1.1500 ;
        RECT 1.1600 1.1500 1.2600 1.3950 ;
        RECT 1.1600 1.3950 1.3300 1.4850 ;
    END
    ANTENNAGATEAREA 0.1272 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6300 0.4900 3.7500 1.7200 ;
    END
    ANTENNADIFFAREA 0.27625 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0050 2.1500 1.3400 ;
        RECT 1.9650 1.3400 2.1500 1.4400 ;
        RECT 1.9650 1.4400 2.0650 1.8150 ;
        RECT 1.9650 1.8150 2.7500 1.9150 ;
        RECT 2.6500 1.4250 2.7500 1.8150 ;
        RECT 2.6500 1.3250 3.0850 1.4250 ;
    END
    ANTENNAGATEAREA 0.1113 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 0.9700 0.7550 1.3700 ;
    END
    ANTENNAGATEAREA 0.0909 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.4300 1.7700 0.5300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6050 0.7600 1.6950 1.6800 ;
      RECT 1.3300 0.6700 1.6950 0.7600 ;
      RECT 2.2150 1.5400 2.3700 1.7100 ;
      RECT 2.2800 0.7800 2.3700 1.5400 ;
      RECT 2.1400 0.6900 2.3700 0.7800 ;
      RECT 2.4700 0.8900 3.1650 0.9800 ;
      RECT 3.0750 0.9800 3.1650 1.1700 ;
      RECT 1.0650 1.9000 1.4450 1.9900 ;
      RECT 1.3550 1.8850 1.4450 1.9000 ;
      RECT 1.3550 1.7950 1.8750 1.8850 ;
      RECT 1.7850 0.5700 1.8750 1.7950 ;
      RECT 1.0350 0.4100 1.4100 0.4800 ;
      RECT 1.3200 0.5000 2.5600 0.5700 ;
      RECT 2.4700 0.5700 2.5600 0.8900 ;
      RECT 1.0350 0.4800 2.5600 0.5000 ;
      RECT 2.4700 0.9800 2.5600 1.6200 ;
      RECT 3.0400 1.6150 3.3500 1.7050 ;
      RECT 3.2600 0.7700 3.3500 1.6150 ;
      RECT 2.9600 0.6800 3.3500 0.7700 ;
      RECT 2.8400 1.8300 3.5300 1.9200 ;
      RECT 2.8400 1.5500 2.9300 1.8300 ;
      RECT 3.4400 0.5700 3.5300 1.8300 ;
      RECT 2.7000 0.4800 3.5300 0.5700 ;
      RECT 2.7000 0.5700 2.8700 0.7900 ;
      RECT 0.0500 1.5100 1.0000 1.6000 ;
      RECT 0.9100 1.2600 1.0000 1.5100 ;
      RECT 0.0500 1.6000 0.1700 1.9600 ;
      RECT 0.0500 0.6300 0.1400 1.5100 ;
      RECT 0.0500 0.5400 0.2450 0.6300 ;
      RECT 0.7150 1.7000 1.2250 1.7900 ;
      RECT 1.1350 1.6850 1.2250 1.7000 ;
      RECT 1.1350 1.5950 1.5100 1.6850 ;
      RECT 1.4200 0.9500 1.5100 1.5950 ;
      RECT 1.1300 0.8600 1.5100 0.9500 ;
      RECT 1.1300 0.6800 1.2200 0.8600 ;
      RECT 0.6350 0.5900 1.2200 0.6800 ;
      RECT 0.7150 1.7900 0.8850 1.9900 ;
  END
END XOR3_X1M_A12TH

MACRO XOR3_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7150 ;
        RECT 0.8550 0.3200 0.9550 0.4950 ;
        RECT 4.7650 0.3200 4.9900 0.3800 ;
        RECT 5.4250 0.3200 5.5250 0.7450 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.8600 1.6550 0.9500 2.0800 ;
        RECT 0.3350 1.6350 0.4350 2.0800 ;
        RECT 5.4250 1.6000 5.5250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0550 1.2500 4.4950 1.3500 ;
        RECT 4.0550 1.1250 4.1550 1.2500 ;
        RECT 3.5500 1.0250 4.1550 1.1250 ;
    END
    ANTENNAGATEAREA 0.1419 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1700 1.2500 5.5500 1.3500 ;
        RECT 5.1700 1.3500 5.2700 1.7950 ;
        RECT 5.4500 0.9450 5.5500 1.2500 ;
        RECT 5.1700 0.8450 5.5500 0.9450 ;
        RECT 5.1700 0.4300 5.2700 0.8450 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8500 1.3050 0.9500 ;
        RECT 1.2050 0.9500 1.3050 1.0400 ;
        RECT 0.2350 0.9500 0.3350 1.1450 ;
        RECT 1.2050 1.0400 1.6050 1.1300 ;
    END
    ANTENNAGATEAREA 0.1716 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.9400 1.1500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.0550 1.2550 1.7900 1.3450 ;
      RECT 1.7000 1.2250 1.7900 1.2550 ;
      RECT 1.7000 1.1350 2.1950 1.2250 ;
      RECT 0.0550 1.3450 0.1700 1.8200 ;
      RECT 0.0550 0.7800 0.1450 1.2550 ;
      RECT 0.0550 0.4100 0.1700 0.7800 ;
      RECT 0.6000 1.4700 2.4600 1.5600 ;
      RECT 2.3700 1.2650 2.4600 1.4700 ;
      RECT 2.3700 1.1750 2.7600 1.2650 ;
      RECT 2.3700 0.9300 2.4600 1.1750 ;
      RECT 1.5750 0.8400 2.4600 0.9300 ;
      RECT 1.5750 0.7500 1.6650 0.8400 ;
      RECT 0.6000 0.6600 1.6650 0.7500 ;
      RECT 0.6000 1.5600 0.6900 1.8750 ;
      RECT 0.6000 0.5000 0.6900 0.6600 ;
      RECT 1.3100 1.6500 2.9600 1.7400 ;
      RECT 2.8700 0.7500 2.9600 1.6500 ;
      RECT 1.8750 0.6600 2.9600 0.7500 ;
      RECT 3.3550 1.2600 3.9450 1.3500 ;
      RECT 3.3550 1.3500 3.4450 1.9450 ;
      RECT 3.3550 0.9050 3.4450 1.2600 ;
      RECT 3.2550 0.8150 3.4450 0.9050 ;
      RECT 3.5850 0.7250 4.3300 0.8150 ;
      RECT 4.2400 0.8150 4.3300 0.8650 ;
      RECT 4.2400 0.8650 4.7200 0.9550 ;
      RECT 4.6300 0.9550 4.7200 1.4400 ;
      RECT 3.9100 1.4400 4.7200 1.5300 ;
      RECT 1.0600 1.8300 3.1400 1.9200 ;
      RECT 3.0500 0.7250 3.1400 1.8300 ;
      RECT 3.0500 0.5700 3.1400 0.6350 ;
      RECT 1.0650 0.4800 3.1400 0.5700 ;
      RECT 3.0500 0.6350 3.6750 0.7250 ;
      RECT 3.9100 1.5300 4.0000 1.7200 ;
      RECT 4.4700 1.6300 4.9000 1.7200 ;
      RECT 4.8100 0.7550 4.9000 1.6300 ;
      RECT 4.4400 0.6650 4.9000 0.7550 ;
      RECT 4.9900 1.0500 5.2700 1.1400 ;
      RECT 3.6300 1.8300 5.0800 1.9200 ;
      RECT 4.1650 1.6300 4.3350 1.8300 ;
      RECT 4.9900 1.1400 5.0800 1.8300 ;
      RECT 4.9900 0.5750 5.0800 1.0500 ;
      RECT 3.8100 0.5250 5.0800 0.5750 ;
      RECT 3.5200 0.4850 5.0800 0.5250 ;
      RECT 3.6300 1.5100 3.7200 1.8300 ;
      RECT 3.5200 0.4350 3.9000 0.4850 ;
  END
END XOR3_X1P4M_A12TH

MACRO XOR3_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7150 ;
        RECT 0.8550 0.3200 0.9550 0.4500 ;
        RECT 5.3150 0.3200 5.4150 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 5.3150 1.7700 5.4150 2.0800 ;
        RECT 0.8600 1.7300 0.9500 2.0800 ;
        RECT 0.3350 1.7000 0.4350 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9000 1.2500 4.3950 1.3500 ;
        RECT 3.9000 1.1250 4.0000 1.2500 ;
        RECT 3.4850 1.0250 4.0000 1.1250 ;
    END
    ANTENNAGATEAREA 0.1689 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0600 1.2500 5.5500 1.3500 ;
        RECT 5.0600 1.3500 5.1600 1.7200 ;
        RECT 5.4500 0.9500 5.5500 1.2500 ;
        RECT 5.0600 0.8500 5.5500 0.9500 ;
        RECT 5.0600 0.4900 5.1600 0.8500 ;
    END
    ANTENNADIFFAREA 0.326 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8500 1.2950 0.9500 ;
        RECT 1.1950 0.9500 1.2950 1.0500 ;
        RECT 0.2350 0.9500 0.3350 1.1450 ;
        RECT 1.1950 1.0500 1.6300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2061 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.0550 1.2550 1.8350 1.3450 ;
      RECT 1.7450 1.2350 1.8350 1.2550 ;
      RECT 1.7450 1.1450 2.1450 1.2350 ;
      RECT 0.0550 1.3450 0.1700 1.7800 ;
      RECT 0.0550 0.7800 0.1450 1.2550 ;
      RECT 0.0550 0.4100 0.1750 0.7800 ;
      RECT 0.6050 1.4450 2.3800 1.5350 ;
      RECT 2.2900 1.1800 2.3800 1.4450 ;
      RECT 2.2900 1.0900 2.6600 1.1800 ;
      RECT 2.2900 0.9300 2.3800 1.0900 ;
      RECT 1.5800 0.8400 2.3800 0.9300 ;
      RECT 1.5800 0.7500 1.6700 0.8400 ;
      RECT 0.6000 0.6600 1.6700 0.7500 ;
      RECT 0.6000 1.6300 0.6900 1.9700 ;
      RECT 0.6000 1.5400 0.6950 1.6300 ;
      RECT 0.6050 1.5350 0.6950 1.5400 ;
      RECT 0.6000 0.5000 0.6900 0.6600 ;
      RECT 1.3100 1.6250 2.8550 1.7150 ;
      RECT 2.7650 0.7500 2.8550 1.6250 ;
      RECT 1.8450 0.6600 2.8550 0.7500 ;
      RECT 3.2250 1.2600 3.7900 1.3500 ;
      RECT 3.2250 1.3500 3.3150 1.8250 ;
      RECT 3.2250 0.7800 3.3150 1.2600 ;
      RECT 3.4650 0.7650 4.2450 0.8550 ;
      RECT 4.1550 0.8550 4.2450 0.9250 ;
      RECT 4.1550 0.9250 4.6100 1.0150 ;
      RECT 4.5200 1.0150 4.6100 1.4400 ;
      RECT 3.7350 1.4400 4.6100 1.5300 ;
      RECT 1.1100 1.8250 3.0350 1.9150 ;
      RECT 1.1100 1.7000 1.2000 1.8250 ;
      RECT 2.9450 0.6900 3.0350 1.8250 ;
      RECT 2.9450 0.5700 3.0350 0.6000 ;
      RECT 1.0650 0.4800 3.0350 0.5700 ;
      RECT 2.9450 0.6000 3.5550 0.6900 ;
      RECT 3.4650 0.6900 3.5550 0.7650 ;
      RECT 3.7350 1.5300 3.8250 1.7200 ;
      RECT 4.3700 1.6300 4.7900 1.7200 ;
      RECT 4.7000 0.7850 4.7900 1.6300 ;
      RECT 4.3750 0.6950 4.7900 0.7850 ;
      RECT 4.8800 1.0500 5.2200 1.1400 ;
      RECT 3.4750 1.8300 4.9700 1.9200 ;
      RECT 4.0550 1.6300 4.2250 1.8300 ;
      RECT 4.8800 1.1400 4.9700 1.8300 ;
      RECT 4.8800 0.5750 4.9700 1.0500 ;
      RECT 3.7100 0.5100 4.9700 0.5750 ;
      RECT 3.4250 0.4850 4.9700 0.5100 ;
      RECT 4.0600 0.4800 4.2300 0.4850 ;
      RECT 3.4750 1.5100 3.5650 1.8300 ;
      RECT 3.4250 0.4200 3.8000 0.4850 ;
  END
END XOR3_X2M_A12TH

MACRO XOR3_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7300 ;
        RECT 0.6050 0.3200 0.7150 0.7400 ;
        RECT 1.1100 0.3200 1.2800 0.5150 ;
        RECT 2.9550 0.3200 3.1250 0.3900 ;
        RECT 3.5200 0.3200 3.6900 0.3900 ;
        RECT 5.4000 0.3200 5.6100 0.3700 ;
        RECT 5.9200 0.3200 6.1300 0.3700 ;
        RECT 6.5100 0.3200 6.6100 0.6650 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 6.5100 1.7700 6.6100 2.0800 ;
        RECT 1.1500 1.7350 1.2400 2.0800 ;
        RECT 0.0900 1.5400 0.1900 2.0800 ;
        RECT 0.6250 1.5100 0.7250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8950 1.0500 4.7950 1.1500 ;
        RECT 4.6950 1.1500 4.7950 1.2600 ;
        RECT 4.6950 1.2600 5.1450 1.3500 ;
    END
    ANTENNAGATEAREA 0.2436 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2550 1.2500 6.9000 1.3500 ;
        RECT 6.2550 1.3500 6.3550 1.7200 ;
        RECT 6.7750 1.3500 6.9000 1.7200 ;
        RECT 6.8000 0.9450 6.9000 1.2500 ;
        RECT 6.2500 0.8450 6.9000 0.9450 ;
        RECT 6.2500 0.5200 6.3500 0.8450 ;
        RECT 6.7750 0.5200 6.9000 0.8450 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7500 1.1500 ;
        RECT 0.6500 0.9500 0.7500 1.0500 ;
        RECT 0.6500 0.8500 1.6650 0.9500 ;
        RECT 1.5650 0.9500 1.6650 1.0200 ;
        RECT 1.5650 1.0200 1.9850 1.1200 ;
    END
    ANTENNAGATEAREA 0.2856 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 1.3650 1.1500 ;
    END
    ANTENNAGATEAREA 0.2205 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.0650 1.2750 2.2700 1.3650 ;
      RECT 2.1800 1.1300 2.2700 1.2750 ;
      RECT 2.1800 1.0400 2.7350 1.1300 ;
      RECT 0.0650 0.9300 0.1550 1.2750 ;
      RECT 0.3550 1.3650 0.4450 1.8700 ;
      RECT 0.0650 0.8400 0.4850 0.9300 ;
      RECT 0.3150 0.4500 0.4850 0.8400 ;
      RECT 0.8900 1.5450 2.0350 1.6250 ;
      RECT 0.8900 1.5350 2.9250 1.5450 ;
      RECT 1.9450 1.4550 2.9250 1.5350 ;
      RECT 2.8350 1.1200 2.9250 1.4550 ;
      RECT 2.8350 1.0300 3.2050 1.1200 ;
      RECT 2.8350 0.9300 2.9250 1.0300 ;
      RECT 1.9500 0.8400 2.9250 0.9300 ;
      RECT 1.9500 0.7500 2.0400 0.8400 ;
      RECT 0.8500 0.6600 2.0400 0.7500 ;
      RECT 1.4100 1.6250 1.5000 1.9450 ;
      RECT 1.3700 0.4600 1.5400 0.6600 ;
      RECT 0.8900 1.6250 0.9800 1.9450 ;
      RECT 0.8500 0.4600 1.0200 0.6600 ;
      RECT 2.1550 1.6500 3.3850 1.7400 ;
      RECT 3.2950 0.7500 3.3850 1.6500 ;
      RECT 2.1600 0.6600 3.3850 0.7500 ;
      RECT 3.8650 1.3500 3.9550 1.7400 ;
      RECT 3.6950 1.2600 4.5600 1.3500 ;
      RECT 3.6950 0.8400 4.0100 0.9300 ;
      RECT 3.6950 0.9300 3.7850 1.2600 ;
      RECT 4.1400 0.8500 5.4200 0.9400 ;
      RECT 5.3300 0.9400 5.4200 1.0800 ;
      RECT 5.3300 1.0800 5.7300 1.1700 ;
      RECT 5.3300 1.1700 5.4200 1.4400 ;
      RECT 4.4150 1.4400 5.4200 1.5300 ;
      RECT 1.6250 1.8300 3.5950 1.9200 ;
      RECT 3.5050 0.7500 3.5950 1.8300 ;
      RECT 3.5050 0.5700 3.5950 0.6600 ;
      RECT 1.6500 0.4800 3.5950 0.5700 ;
      RECT 3.5050 0.6600 4.2300 0.7500 ;
      RECT 4.1400 0.7500 4.2300 0.8500 ;
      RECT 4.4150 1.5300 4.5050 1.6750 ;
      RECT 4.8800 1.6200 5.9350 1.7100 ;
      RECT 5.8450 0.7550 5.9350 1.6200 ;
      RECT 4.3500 0.6650 5.9350 0.7550 ;
      RECT 6.0350 1.0500 6.5850 1.1400 ;
      RECT 4.1550 1.8300 6.1250 1.9200 ;
      RECT 6.0350 1.1400 6.1250 1.8300 ;
      RECT 6.0350 0.5700 6.1250 1.0500 ;
      RECT 4.0950 0.4800 6.1250 0.5700 ;
      RECT 4.1550 1.4900 4.2450 1.8300 ;
  END
END XOR3_X3M_A12TH

MACRO XOR3_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7300 ;
        RECT 0.6050 0.3200 0.7150 0.7200 ;
        RECT 1.1100 0.3200 1.2800 0.5500 ;
        RECT 7.4800 0.3200 7.5800 0.6650 ;
        RECT 8.0000 0.3200 8.1000 0.6650 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 1.1500 1.8100 1.2400 2.0800 ;
        RECT 7.4800 1.7700 7.5800 2.0800 ;
        RECT 8.0000 1.7700 8.1000 2.0800 ;
        RECT 0.0950 1.5800 0.1850 2.0800 ;
        RECT 0.6300 1.5800 0.7200 2.0800 ;
        RECT 4.5500 1.4800 4.7200 2.0800 ;
        RECT 4.0700 1.3850 4.1600 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5300 1.0500 6.1150 1.1500 ;
    END
    ANTENNAGATEAREA 0.2958 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2250 1.2500 7.9500 1.3500 ;
        RECT 7.2250 1.3500 7.3250 1.7200 ;
        RECT 7.7400 1.3500 7.8400 1.7200 ;
        RECT 7.8500 0.9500 7.9500 1.2500 ;
        RECT 7.2200 0.8500 7.9500 0.9500 ;
        RECT 7.2200 0.5000 7.3200 0.8500 ;
        RECT 7.7400 0.5000 7.8400 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7500 1.1500 ;
        RECT 0.6500 0.9500 0.7500 1.0500 ;
        RECT 0.6500 0.8500 1.6650 0.9500 ;
        RECT 1.5650 0.9500 1.6650 1.0500 ;
        RECT 1.5650 1.0500 1.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.3576 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 1.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2736 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.8500 1.6050 2.3400 1.6950 ;
      RECT 2.2500 1.5350 2.3400 1.6050 ;
      RECT 2.2500 1.4450 3.1850 1.5350 ;
      RECT 3.0950 1.1250 3.1850 1.4450 ;
      RECT 3.0950 1.0250 3.6200 1.1250 ;
      RECT 3.0950 0.9500 3.1850 1.0250 ;
      RECT 1.9500 0.8600 3.1850 0.9500 ;
      RECT 1.9500 0.7500 2.0400 0.8600 ;
      RECT 0.8500 0.6600 2.0400 0.7500 ;
      RECT 1.3700 1.6950 1.5400 1.9250 ;
      RECT 1.3700 0.4600 1.5400 0.6600 ;
      RECT 0.8500 1.6950 1.0200 1.9250 ;
      RECT 0.8500 0.4600 1.0200 0.6600 ;
      RECT 2.4500 1.6500 3.8000 1.7400 ;
      RECT 3.7100 0.7500 3.8000 1.6500 ;
      RECT 2.5550 0.6600 3.8000 0.7500 ;
      RECT 4.3300 1.2900 5.5150 1.3800 ;
      RECT 4.3300 1.3800 4.4200 1.7250 ;
      RECT 4.3300 0.6800 4.4200 1.2900 ;
      RECT 1.6500 0.4800 4.6000 0.5700 ;
      RECT 4.5100 0.5700 4.6000 0.8400 ;
      RECT 4.5100 0.8400 6.5950 0.9300 ;
      RECT 6.5050 0.9300 6.5950 1.4150 ;
      RECT 5.6500 1.4150 6.5950 1.5050 ;
      RECT 5.6500 1.5050 5.7400 1.5250 ;
      RECT 4.8700 1.5250 5.7400 1.6150 ;
      RECT 4.8700 1.6150 4.9600 1.9650 ;
      RECT 1.6300 1.8300 3.9800 1.9200 ;
      RECT 3.8900 0.5700 3.9800 1.8300 ;
      RECT 2.2500 0.5700 2.4200 0.7700 ;
      RECT 5.8500 1.6300 6.7950 1.7200 ;
      RECT 6.7050 0.7500 6.7950 1.6300 ;
      RECT 5.0600 0.6600 6.7950 0.7500 ;
      RECT 7.0050 1.0500 7.5400 1.1400 ;
      RECT 5.0650 1.8300 7.0950 1.9200 ;
      RECT 7.0050 1.1400 7.0950 1.8300 ;
      RECT 7.0050 0.5700 7.0950 1.0500 ;
      RECT 4.8300 0.4800 7.0950 0.5700 ;
      RECT 0.0650 1.3900 2.1600 1.4800 ;
      RECT 2.0700 1.1450 2.1600 1.3900 ;
      RECT 2.0700 1.0550 2.8900 1.1450 ;
      RECT 0.0650 0.9300 0.1550 1.3900 ;
      RECT 0.3550 1.4800 0.4450 1.8750 ;
      RECT 0.0650 0.8400 0.4850 0.9300 ;
      RECT 0.3150 0.4500 0.4850 0.8400 ;
  END
END XOR3_X4M_A12TH

MACRO SDFFYQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0700 0.3200 0.1800 0.4250 ;
        RECT 0.9100 0.3200 1.0100 0.6250 ;
        RECT 3.3900 0.3200 3.5600 0.3750 ;
        RECT 4.5850 0.3200 4.7550 0.3600 ;
        RECT 5.1050 0.3200 5.2750 0.3750 ;
        RECT 5.6950 0.3200 5.7950 0.7150 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1950 0.9500 1.3900 ;
        RECT 0.7500 1.0350 0.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.9700 5.1500 1.3000 ;
        RECT 4.3600 1.3000 5.1500 1.4000 ;
        RECT 4.3250 0.8700 5.1500 0.9700 ;
        RECT 4.3600 1.4000 4.4600 1.7100 ;
        RECT 4.8800 1.4000 4.9800 1.7100 ;
        RECT 4.3250 0.6650 4.4950 0.8700 ;
        RECT 4.8450 0.6650 5.0150 0.8700 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 1.0200 5.9600 1.5000 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0500 1.3600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0350 0.3500 1.4600 ;
    END
    ANTENNAGATEAREA 0.0792 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.8750 1.8950 1.0450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.8200 0.7550 1.9200 ;
      RECT 0.4000 0.4200 0.7750 0.5200 ;
      RECT 0.0450 0.5350 0.5000 0.6350 ;
      RECT 0.4000 0.5200 0.5000 0.5350 ;
      RECT 0.0500 1.8000 0.1500 1.8200 ;
      RECT 0.0450 1.6800 0.1500 1.8000 ;
      RECT 0.0450 0.6350 0.1450 1.6800 ;
      RECT 1.3350 1.7300 1.5050 1.9650 ;
      RECT 0.4500 1.6400 1.5050 1.7300 ;
      RECT 0.3650 0.8000 1.4700 0.9000 ;
      RECT 1.3700 0.4800 1.4700 0.8000 ;
      RECT 0.4500 0.9250 0.5400 1.6400 ;
      RECT 0.3650 0.9000 0.5400 0.9250 ;
      RECT 1.6450 1.5450 1.9100 1.6350 ;
      RECT 1.8200 1.0200 1.9100 1.5450 ;
      RECT 1.8200 0.9300 2.4500 1.0200 ;
      RECT 2.3600 1.0200 2.4500 1.2300 ;
      RECT 1.8200 0.8550 1.9100 0.9300 ;
      RECT 1.7400 0.6850 1.9100 0.8550 ;
      RECT 2.0650 1.5450 2.6300 1.6350 ;
      RECT 2.0650 1.1400 2.1550 1.5450 ;
      RECT 2.5400 0.7400 2.6300 1.5450 ;
      RECT 3.5250 1.1200 3.6350 1.3100 ;
      RECT 3.5250 0.9250 3.6150 1.1200 ;
      RECT 2.7250 0.8350 3.6150 0.9250 ;
      RECT 2.7250 0.9250 2.8150 1.7100 ;
      RECT 3.7950 1.0800 4.8300 1.1800 ;
      RECT 3.3100 1.5000 3.8850 1.5900 ;
      RECT 3.7950 1.1800 3.8850 1.5000 ;
      RECT 3.3100 1.0200 3.4000 1.5000 ;
      RECT 3.7950 0.9550 3.8850 1.0800 ;
      RECT 3.7050 0.6650 3.8850 0.9550 ;
      RECT 1.5600 0.4850 5.4850 0.5750 ;
      RECT 5.3950 0.5750 5.4850 1.7100 ;
      RECT 1.5600 1.3250 1.7300 1.4350 ;
      RECT 1.5600 0.5750 1.6500 1.3250 ;
      RECT 3.0550 0.4400 3.2250 0.4850 ;
      RECT 1.7700 1.8300 6.1550 1.9200 ;
      RECT 5.9850 1.6300 6.1550 1.8300 ;
      RECT 6.0650 0.9050 6.1550 1.6300 ;
      RECT 5.5800 0.8150 6.1550 0.9050 ;
      RECT 6.0250 0.5200 6.1550 0.8150 ;
      RECT 5.5800 0.9050 5.6700 1.2400 ;
      RECT 3.0800 1.0250 3.1700 1.8300 ;
  END
END SDFFYQ_X4M_A12TH

MACRO TIEHI_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7200 ;
        RECT 0.6300 0.3200 0.7200 0.7200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 1.3900 0.7500 1.8300 ;
    END
    ANTENNADIFFAREA 0.1456 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3700 1.7600 0.4600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8100 0.1700 1.4700 ;
      RECT 0.4700 0.8900 0.5600 1.2100 ;
      RECT 0.3700 0.8000 0.5600 0.8900 ;
      RECT 0.3700 0.5100 0.4600 0.8000 ;
  END
END TIEHI_X1M_A12TH

MACRO TIELO_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.5850 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6250 0.4400 0.7550 0.9900 ;
    END
    ANTENNADIFFAREA 0.1232 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0800 1.5550 0.1700 2.0800 ;
        RECT 0.6250 1.5550 0.7150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7900 0.1700 1.4650 ;
      RECT 0.3400 1.4800 0.4300 1.7650 ;
      RECT 0.3400 1.3900 0.5600 1.4800 ;
      RECT 0.4700 1.0700 0.5600 1.3900 ;
  END
END TIELO_X1M_A12TH

MACRO WELLANTENNA2_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.4450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.4450 0.3200 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.1500 0.4800 0.2500 1.9200 ;
  END
END WELLANTENNA2_A12TH

MACRO XNOR2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1900 0.8500 1.5500 0.9500 ;
        RECT 1.1900 0.9500 1.2800 1.1600 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2500 1.5150 1.3500 ;
        RECT 0.8500 1.0900 0.9500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7500 0.7500 1.4500 ;
        RECT 0.6500 1.4500 0.8400 1.5500 ;
        RECT 0.6500 0.6600 0.8350 0.7500 ;
    END
    ANTENNADIFFAREA 0.13 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.3700 1.4700 0.5600 1.5600 ;
      RECT 0.4700 0.7500 0.5600 1.4700 ;
      RECT 0.3700 0.6600 0.5600 0.7500 ;
      RECT 0.1700 1.6500 1.1200 1.7400 ;
      RECT 0.9500 1.4400 1.1200 1.6500 ;
      RECT 0.1700 0.4800 1.1100 0.5700 ;
      RECT 0.1700 0.5700 0.2600 1.6500 ;
      RECT 0.5500 1.8300 1.7450 1.9200 ;
      RECT 1.6300 1.4000 1.7450 1.8300 ;
      RECT 1.6550 0.7650 1.7450 1.4000 ;
      RECT 1.6300 0.6650 1.7450 0.7650 ;
      RECT 1.2300 0.5750 1.7450 0.6650 ;
      RECT 1.2300 0.6650 1.3250 0.6700 ;
      RECT 1.0100 0.6700 1.3250 0.7600 ;
      RECT 1.0100 0.7600 1.1000 0.8700 ;
      RECT 0.8400 0.8700 1.1000 0.9600 ;
      RECT 0.5500 1.9200 0.7200 1.9750 ;
  END
END XNOR2_X0P5M_A12TH

MACRO XNOR2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0700 0.3200 0.1700 0.8350 ;
        RECT 1.2550 0.3200 1.4250 0.4900 ;
        RECT 1.5600 0.3200 1.6600 0.4800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7600 0.7500 1.6400 ;
        RECT 0.6500 1.6400 1.0450 1.7400 ;
        RECT 0.6500 0.6600 0.8500 0.7600 ;
    END
    ANTENNADIFFAREA 0.220675 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4300 0.9600 1.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.5450 1.7850 1.6450 2.0800 ;
        RECT 0.0700 1.7550 0.1700 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.0500 1.7500 1.5000 ;
        RECT 1.1250 1.5000 1.7500 1.5900 ;
        RECT 1.1250 1.1700 1.2150 1.5000 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4400 0.6800 0.5300 1.7200 ;
      RECT 1.2050 1.9200 1.3750 1.9900 ;
      RECT 0.2600 1.8300 1.3750 1.9200 ;
      RECT 1.2050 1.7000 1.3750 1.8300 ;
      RECT 0.2600 0.4800 1.0950 0.5700 ;
      RECT 1.0050 0.5700 1.0950 0.7400 ;
      RECT 0.2600 0.5700 0.3500 1.8300 ;
      RECT 1.8300 1.7050 1.9550 1.9600 ;
      RECT 1.8650 0.7000 1.9550 1.7050 ;
      RECT 1.2300 0.6000 1.9550 0.7000 ;
      RECT 1.7850 0.4300 1.9550 0.6000 ;
      RECT 0.8500 1.0300 0.9500 1.5100 ;
      RECT 1.2300 0.7000 1.3300 0.9300 ;
      RECT 0.8500 0.9300 1.3300 1.0300 ;
  END
END XNOR2_X0P7M_A12TH

MACRO XNOR2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0700 0.3200 0.1700 0.6300 ;
        RECT 1.2600 0.3200 1.4300 0.5050 ;
        RECT 1.5600 0.3200 1.6600 0.4450 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7600 0.7500 1.6400 ;
        RECT 0.6500 1.6400 1.0450 1.7400 ;
        RECT 0.6500 0.6600 0.8500 0.7600 ;
    END
    ANTENNADIFFAREA 0.33475 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4300 1.0000 1.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.0200 1.7500 1.5050 ;
        RECT 1.1300 1.5050 1.7500 1.6050 ;
        RECT 1.1300 1.1500 1.2300 1.5050 ;
    END
    ANTENNAGATEAREA 0.1374 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.5450 1.8000 1.6450 2.0800 ;
        RECT 0.0700 1.7700 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4400 0.6800 0.5300 1.7200 ;
      RECT 1.2050 1.9200 1.3750 1.9900 ;
      RECT 0.2600 1.8300 1.3750 1.9200 ;
      RECT 1.2050 1.7000 1.3750 1.8300 ;
      RECT 0.2600 0.4800 1.1650 0.5700 ;
      RECT 0.9950 0.5700 1.1650 0.7100 ;
      RECT 0.9950 0.4200 1.1650 0.4800 ;
      RECT 0.2600 0.5700 0.3500 1.8300 ;
      RECT 1.8250 1.6550 1.9550 1.9000 ;
      RECT 1.8650 0.7200 1.9550 1.6550 ;
      RECT 1.2550 0.6200 1.9550 0.7200 ;
      RECT 1.7950 0.4300 1.9550 0.6200 ;
      RECT 0.8500 0.9500 0.9400 1.5100 ;
      RECT 1.2550 0.7200 1.3550 0.8500 ;
      RECT 0.8500 0.8500 1.3550 0.9500 ;
  END
END XNOR2_X1M_A12TH

MACRO XNOR2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 1.7100 0.3200 1.8000 0.5950 ;
        RECT 2.5100 0.3200 2.6000 0.7600 ;
        RECT 3.0300 0.3200 3.1200 0.8750 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7700 0.7500 1.3750 ;
        RECT 0.6500 1.3750 1.0150 1.4650 ;
        RECT 0.5700 0.5700 0.7500 0.7700 ;
        RECT 0.0900 0.4800 1.2800 0.5700 ;
        RECT 0.0900 0.5700 0.1800 0.8500 ;
    END
    ANTENNADIFFAREA 0.43225 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6350 1.2100 3.0050 1.3500 ;
    END
    ANTENNAGATEAREA 0.1308 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0800 0.3500 1.8200 ;
        RECT 0.2500 1.8200 1.3950 1.9100 ;
        RECT 1.3050 1.9100 1.3950 1.9900 ;
    END
    ANTENNAGATEAREA 0.1854 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.8600 1.7150 1.9500 2.0800 ;
        RECT 2.4400 1.7150 2.5300 2.0800 ;
        RECT 3.0300 1.7150 3.1200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.4800 1.0200 1.5700 1.5500 ;
      RECT 1.0500 0.9550 1.5700 1.0200 ;
      RECT 1.0500 0.9300 1.6000 0.9550 ;
      RECT 1.3900 0.8650 1.6000 0.9300 ;
      RECT 1.6800 1.5150 2.3650 1.6050 ;
      RECT 2.1200 1.6050 2.2100 1.8850 ;
      RECT 2.2750 1.1200 2.3650 1.5150 ;
      RECT 2.1100 1.0300 2.3650 1.1200 ;
      RECT 2.1100 0.6600 2.2000 1.0300 ;
      RECT 0.4700 1.6400 1.7700 1.7300 ;
      RECT 1.6800 1.6050 1.7700 1.6400 ;
      RECT 0.4700 0.9700 0.5600 1.6400 ;
      RECT 0.3500 0.8800 0.5600 0.9700 ;
      RECT 0.3500 0.6600 0.4400 0.8800 ;
      RECT 2.7700 1.5300 2.8600 1.8100 ;
      RECT 2.4550 1.4400 2.8600 1.5300 ;
      RECT 2.3100 0.8500 2.8600 0.9400 ;
      RECT 2.7700 0.5700 2.8600 0.8500 ;
      RECT 2.4550 0.9400 2.5450 1.4400 ;
      RECT 0.8700 0.7750 0.9600 1.1300 ;
      RECT 0.8700 1.1300 1.2200 1.2200 ;
      RECT 1.1300 1.2200 1.2200 1.5500 ;
      RECT 2.3100 0.5700 2.4000 0.8500 ;
      RECT 1.9100 0.4800 2.4000 0.5700 ;
      RECT 1.9100 0.5700 2.0000 0.6850 ;
      RECT 0.8700 0.6850 2.0000 0.7750 ;
      RECT 1.7950 0.7750 1.8850 1.2100 ;
      RECT 1.7950 1.2100 2.1650 1.3000 ;
  END
END XNOR2_X1P4M_A12TH

MACRO XNOR2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.4350 0.3200 0.5350 0.6300 ;
        RECT 0.9700 0.3200 1.0700 0.5800 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.9550 1.8000 1.0550 2.0800 ;
        RECT 0.4350 1.7400 0.5350 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5050 1.0500 0.9950 1.1500 ;
    END
    ANTENNAGATEAREA 0.1872 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 1.7650 1.3500 ;
        RECT 0.2500 1.0550 0.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.252 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.5800 3.3500 1.8200 ;
        RECT 1.1700 1.8200 3.3500 1.9200 ;
        RECT 1.1800 0.4800 3.3500 0.5800 ;
    END
    ANTENNADIFFAREA 0.8515 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0550 0.8550 1.4000 0.9450 ;
      RECT 1.3100 0.9450 1.4000 1.0300 ;
      RECT 1.3100 1.0300 2.0750 1.1200 ;
      RECT 1.9850 1.1200 2.0750 1.2550 ;
      RECT 1.9850 1.2550 2.4400 1.3450 ;
      RECT 0.1150 0.5450 0.2850 0.8550 ;
      RECT 0.1550 1.5650 0.2450 1.8650 ;
      RECT 0.0550 1.4750 0.2450 1.5650 ;
      RECT 0.0550 0.9450 0.1450 1.4750 ;
      RECT 0.7000 1.6100 1.9450 1.7000 ;
      RECT 1.8550 1.5300 1.9450 1.6100 ;
      RECT 1.8550 1.4400 2.8300 1.5300 ;
      RECT 2.7400 0.9400 2.8300 1.4400 ;
      RECT 1.6550 0.8500 2.8300 0.9400 ;
      RECT 1.6550 0.7600 1.7450 0.8500 ;
      RECT 0.6600 0.6700 1.7450 0.7600 ;
      RECT 0.7000 1.7000 0.7900 1.9800 ;
      RECT 0.6600 0.4700 0.8300 0.6700 ;
      RECT 2.0850 1.6400 3.0350 1.7300 ;
      RECT 2.9450 0.7600 3.0350 1.6400 ;
      RECT 2.0300 0.6700 3.0350 0.7600 ;
  END
END XNOR2_X2M_A12TH

MACRO XNOR2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5250 ;
        RECT 0.6150 0.3200 0.7050 0.5250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8050 1.0500 1.2450 1.1500 ;
    END
    ANTENNAGATEAREA 0.2808 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.2900 1.5700 1.3500 ;
        RECT 0.3000 1.2500 1.9400 1.2900 ;
        RECT 1.4700 1.1900 1.9400 1.2500 ;
    END
    ANTENNAGATEAREA 0.3792 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.5700 3.9500 1.8300 ;
        RECT 1.6250 1.8300 3.9500 1.9200 ;
        RECT 1.6300 0.4800 3.9500 0.5700 ;
    END
    ANTENNADIFFAREA 0.8515 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 2.5150 1.6500 3.7250 1.7400 ;
      RECT 3.6350 0.7550 3.7250 1.6500 ;
      RECT 2.4200 0.6650 3.7250 0.7550 ;
      RECT 1.4850 0.9600 2.1200 1.0500 ;
      RECT 2.0300 1.0500 2.1200 1.2100 ;
      RECT 2.0300 1.2100 2.8300 1.3000 ;
      RECT 0.0650 0.8500 1.5750 0.9400 ;
      RECT 1.4850 0.9400 1.5750 0.9600 ;
      RECT 0.0650 0.9400 0.1550 1.5300 ;
      RECT 0.3550 1.6200 0.4450 1.9400 ;
      RECT 0.0650 1.5300 0.4450 1.6200 ;
      RECT 0.3550 0.4400 0.4450 0.8500 ;
      RECT 0.8900 1.4500 3.0700 1.5400 ;
      RECT 1.9050 1.5400 2.0750 1.7400 ;
      RECT 2.9800 1.1200 3.0700 1.4500 ;
      RECT 2.9800 1.0300 3.5250 1.1200 ;
      RECT 2.9800 1.0150 3.0700 1.0300 ;
      RECT 2.2200 0.9250 3.0700 1.0150 ;
      RECT 2.2200 0.7500 2.3100 0.9250 ;
      RECT 0.8500 0.6600 2.3100 0.7500 ;
      RECT 1.4100 1.5400 1.5000 1.8800 ;
      RECT 0.8900 1.5400 0.9800 1.8800 ;
      RECT 0.8500 0.4200 1.0200 0.6600 ;
  END
END XNOR2_X3M_A12TH

MACRO XNOR2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6000 ;
        RECT 0.6100 0.3200 0.7100 0.6000 ;
        RECT 1.1450 0.3200 1.2450 0.5800 ;
        RECT 1.6700 0.3200 1.7600 0.5800 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 1.1450 1.7700 1.2450 2.0800 ;
        RECT 1.6650 1.7700 1.7650 2.0800 ;
        RECT 0.0900 1.7600 0.1900 2.0800 ;
        RECT 0.6100 1.7600 0.7100 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 1.5500 1.1500 ;
    END
    ANTENNAGATEAREA 0.3744 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.2950 2.1500 1.3500 ;
        RECT 0.6500 1.2500 2.6750 1.2950 ;
        RECT 2.0500 1.1950 2.6750 1.2500 ;
        RECT 0.6500 1.1500 0.7500 1.2500 ;
        RECT 0.2600 1.0500 0.7500 1.1500 ;
    END
    ANTENNAGATEAREA 0.498 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 0.5800 5.5500 1.8200 ;
        RECT 1.8750 1.8200 5.5500 1.9200 ;
        RECT 1.8900 0.4800 5.5500 0.5800 ;
        RECT 2.9800 1.6300 3.1500 1.8200 ;
    END
    ANTENNADIFFAREA 1.29675 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 2.7950 1.2500 4.0550 1.3500 ;
      RECT 0.0500 0.8500 2.1500 0.9500 ;
      RECT 2.0500 0.9500 2.1500 0.9550 ;
      RECT 2.0500 0.9550 2.8950 1.0550 ;
      RECT 2.7950 1.0550 2.8950 1.2500 ;
      RECT 0.0500 0.9500 0.1500 1.3100 ;
      RECT 0.3500 1.4100 0.4500 1.7400 ;
      RECT 0.0500 1.3100 0.4500 1.4100 ;
      RECT 0.3500 0.4400 0.4500 0.8500 ;
      RECT 2.7700 1.4450 4.6800 1.5350 ;
      RECT 4.5900 1.1200 4.6800 1.4450 ;
      RECT 4.5900 1.0300 5.0500 1.1200 ;
      RECT 4.5900 1.0150 4.6800 1.0300 ;
      RECT 2.9950 0.9250 4.6800 1.0150 ;
      RECT 2.9950 0.7600 3.0850 0.9250 ;
      RECT 0.8500 0.6700 3.0850 0.7600 ;
      RECT 0.8900 1.5700 2.8600 1.6600 ;
      RECT 2.7700 1.5350 2.8600 1.5700 ;
      RECT 0.8900 1.6600 0.9800 1.9700 ;
      RECT 0.8500 0.4700 1.0200 0.6700 ;
      RECT 1.4100 1.6600 1.5000 1.9600 ;
      RECT 1.3700 0.4700 1.5400 0.6700 ;
      RECT 3.3000 1.6400 5.2600 1.7300 ;
      RECT 5.1700 0.7600 5.2600 1.6400 ;
      RECT 3.1950 0.6700 5.2600 0.7600 ;
  END
END XNOR2_X4M_A12TH

MACRO XNOR3_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 1.8400 1.8300 1.9400 2.0800 ;
        RECT 3.3550 1.8300 3.4650 2.0800 ;
        RECT 0.4000 1.7600 0.4900 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 0.8600 2.1500 1.3500 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6300 0.5750 3.7500 1.9700 ;
    END
    ANTENNADIFFAREA 0.134475 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.2500 1.0000 1.3500 ;
    END
    ANTENNAGATEAREA 0.0453 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.7500 1.5500 ;
        RECT 0.6500 1.5500 0.7500 1.8200 ;
        RECT 0.2500 1.1400 0.3500 1.4500 ;
        RECT 0.6500 1.8200 1.5100 1.9200 ;
        RECT 0.2500 1.0400 0.9600 1.1400 ;
        RECT 1.3400 1.9200 1.5100 1.9850 ;
    END
    ANTENNAGATEAREA 0.0711 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.0500 0.8400 1.1800 0.9300 ;
      RECT 1.0900 0.9300 1.1800 1.0750 ;
      RECT 0.0500 1.6600 0.2450 1.7500 ;
      RECT 0.0500 0.9300 0.1400 1.6600 ;
      RECT 0.0500 0.5550 0.1700 0.8400 ;
      RECT 0.9100 1.5450 1.0000 1.6800 ;
      RECT 0.9100 1.4550 1.4100 1.5450 ;
      RECT 1.3200 0.7500 1.4100 1.4550 ;
      RECT 0.6200 0.6600 1.4100 0.7500 ;
      RECT 1.5000 0.7500 1.5900 1.5300 ;
      RECT 1.5000 0.6600 1.6700 0.7500 ;
      RECT 2.8200 1.9200 2.9900 1.9800 ;
      RECT 2.2400 1.8300 2.9900 1.9200 ;
      RECT 2.2400 0.9600 2.3300 1.8300 ;
      RECT 2.2400 0.8700 2.6350 0.9600 ;
      RECT 2.2400 0.7500 2.3300 0.8700 ;
      RECT 2.0850 0.6600 2.3300 0.7500 ;
      RECT 0.8700 0.4800 2.5300 0.5700 ;
      RECT 2.4400 0.5700 2.5300 0.6800 ;
      RECT 2.4400 0.6800 2.8350 0.7700 ;
      RECT 2.7450 0.7700 2.8350 0.9900 ;
      RECT 2.7450 0.9900 3.1600 1.0800 ;
      RECT 2.7450 1.0800 2.8350 1.4300 ;
      RECT 3.0700 1.0800 3.1600 1.2000 ;
      RECT 2.4900 1.4300 2.8350 1.5200 ;
      RECT 2.4900 1.5200 2.5800 1.6550 ;
      RECT 1.1350 1.6400 1.8750 1.7300 ;
      RECT 1.7850 0.5700 1.8750 1.6400 ;
      RECT 2.9850 1.4600 3.3400 1.5500 ;
      RECT 3.2500 0.7700 3.3400 1.4600 ;
      RECT 2.9450 0.6800 3.3400 0.7700 ;
      RECT 2.7050 1.6400 3.5400 1.7300 ;
      RECT 3.4500 0.5900 3.5400 1.6400 ;
      RECT 2.6550 0.5000 3.5400 0.5900 ;
  END
END XNOR3_X0P5M_A12TH

MACRO XNOR3_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6150 ;
        RECT 3.2300 0.3200 3.4500 0.4100 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.2500 1.0000 1.3500 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0300 0.8500 2.1500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0879 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6300 0.4300 3.7500 1.8300 ;
    END
    ANTENNADIFFAREA 0.187275 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.7500 1.5500 ;
        RECT 0.6500 1.5500 0.7500 1.8200 ;
        RECT 0.2500 1.1400 0.3500 1.4500 ;
        RECT 0.6500 1.8200 1.5100 1.9200 ;
        RECT 0.2500 1.0400 0.9600 1.1400 ;
        RECT 1.3400 1.9200 1.5100 1.9850 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 1.9000 1.8300 1.9900 2.0800 ;
        RECT 3.3250 1.8050 3.4950 2.0800 ;
        RECT 0.4000 1.7100 0.4900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 0.8400 1.1800 0.9300 ;
      RECT 1.0900 0.9300 1.1800 1.1450 ;
      RECT 0.0500 1.6600 0.2450 1.7500 ;
      RECT 0.0500 0.9300 0.1400 1.6600 ;
      RECT 0.0500 0.5050 0.1700 0.8400 ;
      RECT 0.9100 1.5450 1.0000 1.6800 ;
      RECT 0.9100 1.4550 1.4100 1.5450 ;
      RECT 1.3200 0.7500 1.4100 1.4550 ;
      RECT 0.6150 0.6600 1.4100 0.7500 ;
      RECT 1.5000 0.7500 1.5900 1.5300 ;
      RECT 1.5000 0.6600 1.6750 0.7500 ;
      RECT 2.8400 1.9200 3.0100 1.9900 ;
      RECT 2.2600 1.8300 3.0100 1.9200 ;
      RECT 2.2600 0.9700 2.3500 1.8300 ;
      RECT 2.2600 0.8800 2.5150 0.9700 ;
      RECT 2.2600 0.7500 2.3500 0.8800 ;
      RECT 2.0850 0.6600 2.3500 0.7500 ;
      RECT 0.8750 0.4800 2.5300 0.5700 ;
      RECT 2.4400 0.5700 2.5300 0.6800 ;
      RECT 2.4400 0.6800 2.7450 0.7700 ;
      RECT 2.6550 0.7700 2.7450 0.9900 ;
      RECT 2.6550 0.9900 3.1800 1.0800 ;
      RECT 2.6550 1.0800 2.7450 1.3500 ;
      RECT 2.5100 1.3500 2.7450 1.4400 ;
      RECT 2.5100 1.4400 2.6000 1.7400 ;
      RECT 1.1350 1.6400 1.8750 1.7300 ;
      RECT 1.7850 0.5700 1.8750 1.6400 ;
      RECT 3.0200 1.3950 3.3600 1.4850 ;
      RECT 3.2700 0.7750 3.3600 1.3950 ;
      RECT 2.9350 0.6850 3.3600 0.7750 ;
      RECT 2.7150 1.6100 3.5400 1.7000 ;
      RECT 3.4500 0.5900 3.5400 1.6100 ;
      RECT 2.6550 0.5000 3.5400 0.5900 ;
  END
END XNOR3_X0P7M_A12TH

MACRO XNOR3_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4150 0.3200 0.5050 0.6500 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 0.9700 0.7550 1.3700 ;
    END
    ANTENNAGATEAREA 0.0909 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.8900 2.1500 1.4400 ;
    END
    ANTENNAGATEAREA 0.1113 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6300 0.4900 3.7500 1.7200 ;
    END
    ANTENNADIFFAREA 0.27625 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8700 0.3500 1.3600 ;
        RECT 0.2500 0.7700 1.0350 0.8700 ;
        RECT 0.9350 0.8700 1.0350 1.0500 ;
        RECT 0.9350 1.0500 1.2400 1.1500 ;
        RECT 1.1400 1.1500 1.2400 1.3950 ;
        RECT 1.1400 1.3950 1.3300 1.4850 ;
    END
    ANTENNAGATEAREA 0.1272 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.4350 1.7700 0.5250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.5100 1.0000 1.6000 ;
      RECT 0.9100 1.2600 1.0000 1.5100 ;
      RECT 0.0500 1.6000 0.1700 1.9600 ;
      RECT 0.0500 0.6300 0.1400 1.5100 ;
      RECT 0.0500 0.5400 0.2450 0.6300 ;
      RECT 0.7150 1.7000 1.2250 1.7900 ;
      RECT 1.1350 1.6850 1.2250 1.7000 ;
      RECT 1.1350 1.5950 1.5100 1.6850 ;
      RECT 1.4200 0.9500 1.5100 1.5950 ;
      RECT 1.1300 0.8600 1.5100 0.9500 ;
      RECT 1.1300 0.6800 1.2200 0.8600 ;
      RECT 0.6350 0.5900 1.2200 0.6800 ;
      RECT 0.7150 1.7900 0.8850 1.9900 ;
      RECT 1.6050 0.7600 1.6950 1.6800 ;
      RECT 1.3300 0.6700 1.6950 0.7600 ;
      RECT 2.1400 0.6900 2.3700 0.7800 ;
      RECT 2.1600 1.8300 2.7450 1.9200 ;
      RECT 2.2800 0.7800 2.3700 1.6300 ;
      RECT 2.6550 1.4200 2.7450 1.8300 ;
      RECT 2.6550 1.3300 3.0950 1.4200 ;
      RECT 2.1600 1.6300 2.3700 1.9200 ;
      RECT 1.3200 0.5000 2.5600 0.5700 ;
      RECT 2.4700 0.5700 2.5600 0.8900 ;
      RECT 1.0350 0.4800 2.5600 0.5000 ;
      RECT 2.4700 0.8900 3.1650 0.9800 ;
      RECT 2.4700 0.9800 2.5600 1.6200 ;
      RECT 3.0750 0.9800 3.1650 1.1700 ;
      RECT 1.0650 1.9000 1.4450 1.9900 ;
      RECT 1.3550 1.8850 1.4450 1.9000 ;
      RECT 1.3550 1.7950 1.8750 1.8850 ;
      RECT 1.7850 0.5700 1.8750 1.7950 ;
      RECT 1.0350 0.4100 1.4100 0.4800 ;
      RECT 3.0400 1.6150 3.3500 1.7050 ;
      RECT 3.2600 0.7700 3.3500 1.6150 ;
      RECT 2.9600 0.6800 3.3500 0.7700 ;
      RECT 2.8400 1.8300 3.5300 1.9200 ;
      RECT 2.8400 1.5300 2.9300 1.8300 ;
      RECT 3.4400 0.5700 3.5300 1.8300 ;
      RECT 2.7000 0.4800 3.5300 0.5700 ;
      RECT 2.7000 0.5700 2.8700 0.7900 ;
  END
END XNOR3_X1M_A12TH

MACRO XNOR3_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7150 ;
        RECT 0.8550 0.3200 0.9550 0.4950 ;
        RECT 4.7450 0.3200 4.9150 0.3550 ;
        RECT 5.4250 0.3200 5.5250 0.7450 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.9400 1.1500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8500 1.5750 0.9500 ;
        RECT 1.4750 0.9500 1.5750 1.0300 ;
        RECT 0.2350 0.9500 0.3350 1.1450 ;
        RECT 1.4750 1.0300 1.8400 1.1300 ;
        RECT 1.7400 1.1300 1.8400 1.2900 ;
        RECT 1.7400 1.2900 2.1450 1.3800 ;
    END
    ANTENNAGATEAREA 0.1725 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1700 1.2500 5.5500 1.3500 ;
        RECT 5.1700 1.3500 5.2700 1.7950 ;
        RECT 5.4500 0.9450 5.5500 1.2500 ;
        RECT 5.1700 0.8450 5.5500 0.9450 ;
        RECT 5.1700 0.4300 5.2700 0.8450 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.2500 3.9100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1419 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.8600 1.6550 0.9500 2.0800 ;
        RECT 0.3350 1.6350 0.4350 2.0800 ;
        RECT 5.4300 1.6000 5.5200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.2550 1.6050 1.3450 ;
      RECT 0.0550 1.3450 0.1700 1.8200 ;
      RECT 0.0550 0.7800 0.1450 1.2550 ;
      RECT 0.0550 0.4100 0.1700 0.7800 ;
      RECT 0.6000 1.4700 2.4600 1.5600 ;
      RECT 2.3700 1.2650 2.4600 1.4700 ;
      RECT 2.3700 1.1750 2.7600 1.2650 ;
      RECT 2.3700 0.9300 2.4600 1.1750 ;
      RECT 1.7250 0.8400 2.4600 0.9300 ;
      RECT 1.7250 0.7500 1.8150 0.8400 ;
      RECT 0.6000 0.6600 1.8150 0.7500 ;
      RECT 1.3600 1.5600 1.4700 1.7200 ;
      RECT 0.6000 1.5600 0.6900 1.8750 ;
      RECT 0.6000 0.5000 0.6900 0.6600 ;
      RECT 1.8300 1.6500 2.9600 1.7400 ;
      RECT 2.8700 0.7500 2.9600 1.6500 ;
      RECT 1.9250 0.6600 2.9600 0.7500 ;
      RECT 3.2300 1.0300 4.1700 1.1200 ;
      RECT 4.0800 1.1200 4.1700 1.2600 ;
      RECT 4.0800 1.2600 4.4950 1.3500 ;
      RECT 3.3550 1.6250 3.4450 1.9500 ;
      RECT 3.2300 1.5350 3.4450 1.6250 ;
      RECT 3.2300 1.1200 3.3200 1.5350 ;
      RECT 3.2300 0.9050 3.3200 1.0300 ;
      RECT 3.2300 0.8150 3.4450 0.9050 ;
      RECT 3.0500 0.6350 3.6750 0.7250 ;
      RECT 3.5850 0.7250 4.3300 0.8150 ;
      RECT 4.2400 0.8150 4.3300 0.8650 ;
      RECT 4.2400 0.8650 4.7200 0.9550 ;
      RECT 4.6300 0.9550 4.7200 1.4400 ;
      RECT 3.9100 1.4400 4.7200 1.5300 ;
      RECT 3.9100 1.5300 4.0000 1.7200 ;
      RECT 1.0600 1.8300 3.1400 1.9200 ;
      RECT 3.0500 0.7250 3.1400 1.8300 ;
      RECT 3.0500 0.5700 3.1400 0.6350 ;
      RECT 1.0650 0.4800 3.1400 0.5700 ;
      RECT 4.4700 1.6300 4.9000 1.7200 ;
      RECT 4.8100 0.7550 4.9000 1.6300 ;
      RECT 4.4400 0.6650 4.9000 0.7550 ;
      RECT 4.9900 1.0500 5.3300 1.1400 ;
      RECT 3.6300 1.8300 5.0800 1.9200 ;
      RECT 4.1650 1.6300 4.3350 1.8300 ;
      RECT 3.6300 1.5100 3.7200 1.8300 ;
      RECT 4.9900 1.1400 5.0800 1.8300 ;
      RECT 4.9900 0.5700 5.0800 1.0500 ;
      RECT 3.8050 0.5450 5.0800 0.5700 ;
      RECT 3.5400 0.4800 5.0800 0.5450 ;
      RECT 3.5400 0.4550 3.9150 0.4800 ;
  END
END XNOR3_X1P4M_A12TH

MACRO XNOR3_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7150 ;
        RECT 0.8550 0.3200 0.9550 0.4500 ;
        RECT 5.4300 0.3200 5.5200 0.6300 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8500 1.2950 0.9150 ;
        RECT 0.2350 0.9150 1.6450 0.9500 ;
        RECT 0.2350 0.9500 0.3350 1.1450 ;
        RECT 1.1950 0.9500 1.6450 1.0150 ;
    END
    ANTENNAGATEAREA 0.2061 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1700 1.2500 5.5500 1.3500 ;
        RECT 5.1700 1.3500 5.2700 1.7200 ;
        RECT 5.4500 0.9500 5.5500 1.2500 ;
        RECT 5.1700 0.8500 5.5500 0.9500 ;
        RECT 5.1700 0.4900 5.2600 0.8500 ;
    END
    ANTENNADIFFAREA 0.326 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5250 1.2500 3.9450 1.3500 ;
    END
    ANTENNAGATEAREA 0.1689 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 5.4300 1.7700 5.5200 2.0800 ;
        RECT 0.8600 1.7300 0.9500 2.0800 ;
        RECT 0.3350 1.7000 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.2550 1.9550 1.3450 ;
      RECT 1.8650 1.1100 1.9550 1.2550 ;
      RECT 1.8650 1.0200 2.2550 1.1100 ;
      RECT 0.0550 1.3450 0.1700 1.7600 ;
      RECT 0.0550 0.7800 0.1450 1.2550 ;
      RECT 0.0550 0.4100 0.1750 0.7800 ;
      RECT 0.6000 1.5400 1.6600 1.6300 ;
      RECT 1.5700 1.5350 1.6600 1.5400 ;
      RECT 1.5700 1.4450 2.4900 1.5350 ;
      RECT 2.4000 1.1800 2.4900 1.4450 ;
      RECT 2.4000 1.0900 2.7700 1.1800 ;
      RECT 2.4000 0.9300 2.4900 1.0900 ;
      RECT 1.7550 0.8400 2.4900 0.9300 ;
      RECT 1.7550 0.7500 1.8450 0.8400 ;
      RECT 0.6000 0.6600 1.8450 0.7500 ;
      RECT 0.6000 1.6300 0.6900 1.9700 ;
      RECT 0.6000 0.5000 0.6900 0.6600 ;
      RECT 1.8300 1.6250 2.9650 1.7150 ;
      RECT 2.8750 0.7500 2.9650 1.6250 ;
      RECT 1.9550 0.6600 2.9650 0.7500 ;
      RECT 3.2500 1.0150 4.1750 1.1150 ;
      RECT 4.0750 1.1150 4.1750 1.2500 ;
      RECT 4.0750 1.2500 4.5050 1.3500 ;
      RECT 3.3350 1.5900 3.4250 1.9100 ;
      RECT 3.2500 1.5000 3.4250 1.5900 ;
      RECT 3.2500 1.1150 3.3400 1.5000 ;
      RECT 3.2500 0.9150 3.3400 1.0150 ;
      RECT 3.2500 0.8250 3.4650 0.9150 ;
      RECT 3.0550 0.6450 3.6650 0.7350 ;
      RECT 3.5750 0.7350 3.6650 0.7650 ;
      RECT 3.5750 0.7650 4.3550 0.8550 ;
      RECT 4.2650 0.8550 4.3550 0.9250 ;
      RECT 4.2650 0.9250 4.7200 1.0150 ;
      RECT 4.6300 1.0150 4.7200 1.4400 ;
      RECT 3.8450 1.4400 4.7200 1.5300 ;
      RECT 3.8450 1.5300 3.9350 1.7200 ;
      RECT 1.0600 1.8050 3.1450 1.8950 ;
      RECT 3.0550 0.7350 3.1450 1.8050 ;
      RECT 3.0550 0.5700 3.1450 0.6450 ;
      RECT 1.0650 0.4800 3.1450 0.5700 ;
      RECT 4.4800 1.6300 4.9000 1.7200 ;
      RECT 4.8100 0.7850 4.9000 1.6300 ;
      RECT 4.4850 0.6950 4.9000 0.7850 ;
      RECT 4.9900 1.0500 5.3300 1.1400 ;
      RECT 3.5850 1.8300 5.0800 1.9200 ;
      RECT 4.1650 1.6300 4.3350 1.8300 ;
      RECT 3.5850 1.5100 3.6750 1.8300 ;
      RECT 4.9900 1.1400 5.0800 1.8300 ;
      RECT 4.9900 0.5750 5.0800 1.0500 ;
      RECT 3.8450 0.5300 5.0800 0.5750 ;
      RECT 3.5600 0.4850 5.0800 0.5300 ;
      RECT 3.5600 0.4400 3.9350 0.4850 ;
  END
END XNOR3_X2M_A12TH

MACRO XNOR3_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7300 ;
        RECT 0.6050 0.3200 0.7150 0.7400 ;
        RECT 1.1100 0.3200 1.2800 0.5150 ;
        RECT 3.2050 0.3200 3.3750 0.3900 ;
        RECT 3.7700 0.3200 3.9400 0.3900 ;
        RECT 5.6500 0.3200 5.8600 0.3700 ;
        RECT 6.1700 0.3200 6.3800 0.3700 ;
        RECT 6.7600 0.3200 6.8600 0.6650 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 1.3650 1.1500 ;
    END
    ANTENNAGATEAREA 0.2241 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7500 1.1500 ;
        RECT 0.6500 0.9500 0.7500 1.0500 ;
        RECT 0.6500 0.8500 1.6650 0.9500 ;
        RECT 1.5650 0.9500 1.6650 1.0200 ;
        RECT 1.5650 1.0200 1.9650 1.1200 ;
    END
    ANTENNAGATEAREA 0.2868 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5050 1.2500 7.1500 1.3500 ;
        RECT 6.5050 1.3500 6.6050 1.7200 ;
        RECT 7.0250 1.3500 7.1500 1.7200 ;
        RECT 7.0500 0.9450 7.1500 1.2500 ;
        RECT 6.5000 0.8450 7.1500 0.9450 ;
        RECT 6.5000 0.5200 6.6000 0.8450 ;
        RECT 7.0250 0.5200 7.1500 0.8450 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 6.7600 1.7700 6.8600 2.0800 ;
        RECT 1.1500 1.7300 1.2400 2.0800 ;
        RECT 0.0900 1.5400 0.1900 2.0800 ;
        RECT 0.6250 1.5100 0.7250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1600 1.0500 4.7350 1.1500 ;
    END
    ANTENNAGATEAREA 0.2442 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0650 1.2750 2.1450 1.3650 ;
      RECT 2.0550 1.1300 2.1450 1.2750 ;
      RECT 2.0550 1.0400 2.7350 1.1300 ;
      RECT 0.0650 0.9300 0.1550 1.2750 ;
      RECT 0.3550 1.3650 0.4450 1.8700 ;
      RECT 0.0650 0.8400 0.4850 0.9300 ;
      RECT 0.3150 0.4500 0.4850 0.8400 ;
      RECT 0.8900 1.5350 2.2800 1.6200 ;
      RECT 0.8900 1.5300 3.0700 1.5350 ;
      RECT 2.1900 1.4450 3.0700 1.5300 ;
      RECT 2.9800 1.1200 3.0700 1.4450 ;
      RECT 2.9800 1.0300 3.4300 1.1200 ;
      RECT 2.9800 0.9350 3.0700 1.0300 ;
      RECT 2.1550 0.8450 3.0700 0.9350 ;
      RECT 2.1550 0.7500 2.2450 0.8450 ;
      RECT 0.8500 0.6600 2.2450 0.7500 ;
      RECT 1.4100 1.6200 1.5000 1.9400 ;
      RECT 1.3700 0.4600 1.5400 0.6600 ;
      RECT 0.8900 1.6200 0.9800 1.9400 ;
      RECT 0.8500 0.4600 1.0200 0.6600 ;
      RECT 2.3950 1.6500 3.6350 1.7400 ;
      RECT 3.5450 0.7500 3.6350 1.6500 ;
      RECT 2.4000 0.6600 3.6350 0.7500 ;
      RECT 4.1150 1.3500 4.2050 1.7400 ;
      RECT 3.9450 1.2600 5.4300 1.3500 ;
      RECT 3.9450 0.8400 4.2450 0.9300 ;
      RECT 3.9450 0.9300 4.0350 1.2600 ;
      RECT 3.7550 0.6600 4.4800 0.7500 ;
      RECT 4.3900 0.7500 4.4800 0.8500 ;
      RECT 4.3900 0.8500 5.6700 0.9400 ;
      RECT 5.5800 0.9400 5.6700 1.0800 ;
      RECT 5.5800 1.0800 5.9800 1.1700 ;
      RECT 5.5800 1.1700 5.6700 1.4400 ;
      RECT 4.6650 1.4400 5.6700 1.5300 ;
      RECT 4.6650 1.5300 4.7550 1.6750 ;
      RECT 1.6250 1.8300 3.8450 1.9200 ;
      RECT 3.7550 0.7500 3.8450 1.8300 ;
      RECT 3.7550 0.5700 3.8450 0.6600 ;
      RECT 1.6500 0.4800 3.8450 0.5700 ;
      RECT 5.1300 1.6200 6.1850 1.7100 ;
      RECT 6.0950 0.7550 6.1850 1.6200 ;
      RECT 4.6000 0.6650 6.1850 0.7550 ;
      RECT 6.2850 1.0500 6.8350 1.1400 ;
      RECT 4.4050 1.8300 6.3750 1.9200 ;
      RECT 4.4050 1.4900 4.4950 1.8300 ;
      RECT 6.2850 1.1400 6.3750 1.8300 ;
      RECT 6.2850 0.5700 6.3750 1.0500 ;
      RECT 4.3450 0.4800 6.3750 0.5700 ;
  END
END XNOR3_X3M_A12TH

MACRO XNOR3_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7450 ;
        RECT 0.6150 0.3200 0.7050 0.7200 ;
        RECT 1.1100 0.3200 1.2800 0.5500 ;
        RECT 6.3850 0.3200 6.5950 0.3700 ;
        RECT 6.9050 0.3200 7.1150 0.3700 ;
        RECT 7.4850 0.3200 7.5750 0.6650 ;
        RECT 8.0050 0.3200 8.0950 0.6650 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 1.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2736 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7500 1.1500 ;
        RECT 0.6500 0.9500 0.7500 1.0500 ;
        RECT 0.6500 0.8500 1.6650 0.9500 ;
        RECT 1.5650 0.9500 1.6650 1.0650 ;
        RECT 1.5650 1.0650 1.9650 1.1650 ;
    END
    ANTENNAGATEAREA 0.3576 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2250 1.2500 7.9500 1.3500 ;
        RECT 7.2250 1.3500 7.3250 1.7200 ;
        RECT 7.7450 1.3500 7.8350 1.7200 ;
        RECT 7.8500 0.9500 7.9500 1.2500 ;
        RECT 7.2250 0.8500 7.9500 0.9500 ;
        RECT 7.2250 0.5200 7.3150 0.8500 ;
        RECT 7.7450 0.5200 7.8350 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6100 1.0500 5.0400 1.1500 ;
    END
    ANTENNAGATEAREA 0.2958 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 1.1500 1.8100 1.2400 2.0800 ;
        RECT 7.4800 1.7700 7.5800 2.0800 ;
        RECT 8.0000 1.7700 8.1000 2.0800 ;
        RECT 0.0950 1.5800 0.1850 2.0800 ;
        RECT 0.6300 1.5800 0.7200 2.0800 ;
        RECT 4.5500 1.4800 4.7200 2.0800 ;
        RECT 4.0700 1.3900 4.1600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0650 1.3900 2.1550 1.4800 ;
      RECT 2.0650 1.1450 2.1550 1.3900 ;
      RECT 2.0650 1.0550 2.8900 1.1450 ;
      RECT 0.0650 0.9300 0.1550 1.3900 ;
      RECT 0.3550 1.4800 0.4450 1.8700 ;
      RECT 0.0650 0.8400 0.4450 0.9300 ;
      RECT 0.3550 0.4250 0.4450 0.8400 ;
      RECT 0.8500 1.6050 2.3350 1.6950 ;
      RECT 2.2450 1.5350 2.3350 1.6050 ;
      RECT 2.2450 1.4450 3.1850 1.5350 ;
      RECT 3.0950 1.1250 3.1850 1.4450 ;
      RECT 3.0950 1.0250 3.6200 1.1250 ;
      RECT 3.0950 0.9500 3.1850 1.0250 ;
      RECT 1.9500 0.8600 3.1850 0.9500 ;
      RECT 1.9500 0.7500 2.0400 0.8600 ;
      RECT 0.8500 0.6600 2.0400 0.7500 ;
      RECT 1.3700 1.6950 1.5400 1.9100 ;
      RECT 1.3700 0.4600 1.5400 0.6600 ;
      RECT 0.8500 1.6950 1.0200 1.9100 ;
      RECT 0.8500 0.4600 1.0200 0.6600 ;
      RECT 2.4500 1.6500 3.8000 1.7400 ;
      RECT 3.7100 0.7500 3.8000 1.6500 ;
      RECT 2.5550 0.6600 3.8000 0.7500 ;
      RECT 4.3300 1.2900 5.5300 1.3800 ;
      RECT 5.4400 1.1550 5.5300 1.2900 ;
      RECT 5.4400 1.0650 6.1150 1.1550 ;
      RECT 4.3300 1.3800 4.4200 1.7200 ;
      RECT 4.3300 0.6800 4.4200 1.2900 ;
      RECT 4.5100 0.8400 6.5950 0.9300 ;
      RECT 6.5050 0.9300 6.5950 1.4150 ;
      RECT 5.6500 1.4150 6.5950 1.5050 ;
      RECT 5.6500 1.5050 5.7400 1.5250 ;
      RECT 4.8700 1.5250 5.7400 1.6150 ;
      RECT 4.8700 1.6150 4.9600 1.9650 ;
      RECT 1.6500 0.4800 4.6000 0.5700 ;
      RECT 4.5100 0.5700 4.6000 0.8400 ;
      RECT 1.6300 1.8300 3.9800 1.9200 ;
      RECT 3.8900 0.5700 3.9800 1.8300 ;
      RECT 2.2500 0.5700 2.4200 0.7700 ;
      RECT 5.8500 1.6300 6.7950 1.7200 ;
      RECT 6.7050 0.7500 6.7950 1.6300 ;
      RECT 5.0600 0.6600 6.7950 0.7500 ;
      RECT 7.0050 1.0500 7.5400 1.1400 ;
      RECT 5.0650 1.8300 7.0950 1.9200 ;
      RECT 7.0050 1.1400 7.0950 1.8300 ;
      RECT 7.0050 0.5700 7.0950 1.0500 ;
      RECT 4.8300 0.4800 7.0950 0.5700 ;
  END
END XNOR3_X4M_A12TH

MACRO XOR2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 1.2650 0.3200 1.3650 0.5750 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7350 0.8600 1.5600 0.9600 ;
        RECT 0.7350 0.9600 0.8350 1.5200 ;
        RECT 1.0100 0.8500 1.5600 0.8600 ;
        RECT 1.4500 0.7000 1.5600 0.8500 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.0500 1.4300 1.1500 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.3500 1.5300 1.4500 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2100 0.6450 1.3900 ;
        RECT 0.5450 1.3900 0.6450 1.6400 ;
        RECT 0.5450 0.7500 0.6450 1.2100 ;
        RECT 0.5450 1.6400 0.9500 1.7400 ;
        RECT 0.5450 0.6600 0.7700 0.7500 ;
    END
    ANTENNADIFFAREA 0.144625 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2550 1.5400 0.4550 1.7100 ;
      RECT 0.2550 0.6800 0.4550 0.8600 ;
      RECT 0.2550 0.8600 0.3450 1.5400 ;
      RECT 0.0700 1.8300 1.1800 1.9200 ;
      RECT 1.0900 1.5300 1.1800 1.8300 ;
      RECT 0.0700 0.4800 1.0150 0.5700 ;
      RECT 0.9150 0.5700 1.0150 0.7350 ;
      RECT 0.0700 0.5700 0.1600 1.8300 ;
      RECT 1.6300 1.3600 1.7500 1.9300 ;
      RECT 0.9550 1.2700 1.7500 1.3600 ;
      RECT 1.6600 0.5900 1.7500 1.2700 ;
      RECT 1.5650 0.5000 1.7500 0.5900 ;
  END
END XOR2_X0P5M_A12TH

MACRO XOR2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0700 0.3200 0.1700 0.8350 ;
        RECT 1.2900 0.3200 1.3900 0.5400 ;
        RECT 1.5600 0.3200 1.6600 0.4500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7600 0.7500 1.6400 ;
        RECT 0.6500 1.6400 1.0450 1.7400 ;
        RECT 0.6500 0.6600 0.8500 0.7600 ;
    END
    ANTENNADIFFAREA 0.238875 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8500 1.3300 0.9500 ;
        RECT 0.8500 0.9500 0.9500 1.5100 ;
        RECT 1.2300 0.7500 1.3300 0.8500 ;
        RECT 1.2300 0.6500 1.7550 0.7500 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.5450 1.7850 1.6450 2.0800 ;
        RECT 0.0700 1.7550 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4400 0.6800 0.5300 1.7200 ;
      RECT 1.2150 1.9200 1.3850 1.9900 ;
      RECT 0.2600 1.8300 1.3850 1.9200 ;
      RECT 1.2150 1.7000 1.3850 1.8300 ;
      RECT 0.2600 0.5700 0.3500 1.8300 ;
      RECT 0.2600 0.4800 1.1850 0.5700 ;
      RECT 1.8300 1.6000 1.9550 1.9800 ;
      RECT 1.1350 1.5100 1.9550 1.6000 ;
      RECT 1.8650 0.5300 1.9550 1.5100 ;
      RECT 1.7700 0.4400 1.9550 0.5300 ;
      RECT 1.1350 1.1700 1.2250 1.5100 ;
  END
END XOR2_X0P7M_A12TH

MACRO XOR2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0700 0.3200 0.1700 0.6300 ;
        RECT 1.2950 0.3200 1.3950 0.5600 ;
        RECT 1.5600 0.3200 1.6600 0.5600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7600 0.7500 1.6400 ;
        RECT 0.6500 1.6400 1.0450 1.7400 ;
        RECT 0.6500 0.6600 0.8500 0.7600 ;
    END
    ANTENNADIFFAREA 0.34125 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9600 1.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8500 1.3550 0.9500 ;
        RECT 0.8500 0.9500 0.9500 1.5100 ;
        RECT 1.2550 0.7500 1.3550 0.8500 ;
        RECT 1.2550 0.6500 1.7600 0.7500 ;
        RECT 1.6500 0.7500 1.7600 0.9000 ;
    END
    ANTENNAGATEAREA 0.1374 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.5450 1.8000 1.6450 2.0800 ;
        RECT 0.0700 1.7700 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4400 0.6800 0.5300 1.7200 ;
      RECT 1.2150 1.9200 1.3850 1.9900 ;
      RECT 0.2600 1.8300 1.3850 1.9200 ;
      RECT 1.2150 1.7000 1.3850 1.8300 ;
      RECT 0.2600 0.5700 0.3500 1.8300 ;
      RECT 0.2600 0.4800 1.1650 0.5700 ;
      RECT 0.9950 0.5700 1.1650 0.7100 ;
      RECT 0.9950 0.4200 1.1650 0.4800 ;
      RECT 1.8300 1.6000 1.9550 1.9000 ;
      RECT 1.1400 1.5100 1.9550 1.6000 ;
      RECT 1.8650 0.5500 1.9550 1.5100 ;
      RECT 1.7700 0.4600 1.9550 0.5500 ;
      RECT 1.1400 1.1500 1.2300 1.5100 ;
  END
END XOR2_X1M_A12TH

MACRO XOR2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 1.7650 0.3200 1.9750 0.3900 ;
        RECT 2.5100 0.3200 2.6000 0.5750 ;
        RECT 3.0300 0.3200 3.1200 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5250 0.8500 1.2100 0.9500 ;
        RECT 0.5250 0.9500 0.6150 1.2400 ;
        RECT 0.5250 0.7700 0.6900 0.8500 ;
        RECT 1.1200 0.6600 1.2100 0.8500 ;
        RECT 0.5250 1.2400 1.1300 1.3300 ;
        RECT 0.6000 0.5700 0.6900 0.7700 ;
        RECT 1.0400 1.3300 1.1300 1.5300 ;
        RECT 0.0800 0.4800 0.6900 0.5700 ;
        RECT 0.0800 0.5700 0.1700 0.8500 ;
    END
    ANTENNADIFFAREA 0.5278 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7150 1.0500 3.1350 1.1500 ;
    END
    ANTENNAGATEAREA 0.1308 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.9700 2.0100 2.0600 2.0800 ;
        RECT 2.4900 1.8400 2.5800 2.0800 ;
        RECT 3.0100 1.8400 3.1000 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7250 1.0500 1.1900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1854 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.8600 1.6500 1.8600 1.7400 ;
      RECT 1.2400 1.3300 1.3300 1.6500 ;
      RECT 1.2400 1.2400 1.5500 1.3300 ;
      RECT 1.4600 1.1500 1.5500 1.2400 ;
      RECT 1.4600 1.0600 1.6550 1.1500 ;
      RECT 1.5650 0.6600 1.6550 1.0600 ;
      RECT 0.3450 1.1400 0.4350 1.4200 ;
      RECT 0.8600 1.5100 0.9500 1.6500 ;
      RECT 0.3450 1.4200 0.9500 1.5100 ;
      RECT 0.6000 1.8300 2.3600 1.9200 ;
      RECT 2.1800 1.7100 2.3600 1.8300 ;
      RECT 2.1800 1.6200 2.4450 1.7100 ;
      RECT 2.3550 0.9800 2.4450 1.6200 ;
      RECT 2.1100 0.8900 2.4450 0.9800 ;
      RECT 2.1100 0.6600 2.2000 0.8900 ;
      RECT 0.1500 1.0300 0.2400 1.6300 ;
      RECT 0.1500 0.9400 0.4300 1.0300 ;
      RECT 0.3400 0.6600 0.4300 0.9400 ;
      RECT 0.6000 1.7200 0.7700 1.8300 ;
      RECT 0.1500 1.6300 0.7700 1.7200 ;
      RECT 2.7500 1.5400 2.8400 1.9100 ;
      RECT 2.5350 1.4500 2.8400 1.5400 ;
      RECT 2.3100 0.7100 2.8600 0.8000 ;
      RECT 2.7700 0.4300 2.8600 0.7100 ;
      RECT 2.5350 0.8000 2.6250 1.4500 ;
      RECT 2.3100 0.5700 2.4000 0.7100 ;
      RECT 0.8600 0.4800 2.4000 0.5700 ;
      RECT 1.8750 0.5700 1.9650 1.0700 ;
      RECT 1.8750 1.0700 2.2450 1.1600 ;
      RECT 1.8750 1.1600 1.9650 1.4200 ;
      RECT 1.4200 1.4200 1.9650 1.5100 ;
      RECT 1.4200 1.5100 1.6100 1.5600 ;
      RECT 0.8600 0.5700 0.9500 0.7000 ;
  END
END XOR2_X1P4M_A12TH

MACRO XOR2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 1.9100 0.3200 2.0000 0.6000 ;
        RECT 2.4900 0.3200 2.5800 0.6550 ;
        RECT 3.0100 0.3200 3.1000 0.6550 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.0500 1.9000 1.1400 ;
        RECT 0.2550 1.1400 0.6250 1.1650 ;
        RECT 1.8100 1.1400 1.9000 1.2200 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 1.3450 1.5500 ;
        RECT 0.1300 1.5500 0.2200 1.8200 ;
        RECT 0.0750 0.9400 0.1650 1.4500 ;
        RECT 0.0750 0.8500 0.2200 0.9400 ;
        RECT 0.1250 0.5700 0.2200 0.8500 ;
        RECT 0.1250 0.4900 1.2600 0.5700 ;
        RECT 0.6500 0.5700 1.2600 0.5800 ;
        RECT 0.1250 0.4800 0.7400 0.4900 ;
        RECT 1.1700 0.4100 1.2600 0.4900 ;
        RECT 0.6500 0.5800 0.7400 0.7800 ;
        RECT 0.6500 0.4100 0.7400 0.4800 ;
    END
    ANTENNADIFFAREA 0.703125 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.9250 2.0100 2.0150 2.0800 ;
        RECT 2.4900 1.8300 2.5800 2.0800 ;
        RECT 3.0100 1.8300 3.1000 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6100 1.0500 3.0300 1.1500 ;
    END
    ANTENNAGATEAREA 0.183 ;
  END B
  OBS
    LAYER M1 ;
      RECT 1.6300 1.3400 1.7200 1.5600 ;
      RECT 0.8500 1.2500 1.7200 1.3400 ;
      RECT 1.4000 0.5000 1.4900 0.6000 ;
      RECT 1.4000 0.4100 1.7800 0.5000 ;
      RECT 0.8700 1.6500 1.9200 1.7400 ;
      RECT 1.8300 1.4000 1.9200 1.6500 ;
      RECT 1.8300 1.3100 2.1400 1.4000 ;
      RECT 2.0500 0.9600 2.1400 1.3100 ;
      RECT 0.3900 0.8700 2.1400 0.9600 ;
      RECT 0.3900 0.6600 0.4800 0.8700 ;
      RECT 0.3300 1.8300 2.3200 1.9200 ;
      RECT 2.2300 0.7800 2.3200 1.8300 ;
      RECT 0.8500 0.6900 2.3200 0.7800 ;
      RECT 2.2300 0.4100 2.3200 0.6900 ;
      RECT 2.7500 1.3300 2.8400 1.6350 ;
      RECT 2.4100 1.2400 2.8400 1.3300 ;
      RECT 2.4100 0.8700 2.8400 0.9600 ;
      RECT 2.7500 0.5750 2.8400 0.8700 ;
      RECT 2.4100 0.9600 2.5000 1.2400 ;
  END
END XOR2_X2M_A12TH

MACRO XOR2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5600 ;
        RECT 0.6100 0.3200 0.7100 0.7400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.0900 1.8000 0.1900 2.0800 ;
        RECT 0.6100 1.8000 0.7100 2.0800 ;
        RECT 1.1450 1.8000 1.2450 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.3050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2808 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8500 1.6350 0.9500 ;
        RECT 1.5350 0.9500 1.6350 0.9550 ;
        RECT 0.4500 0.9500 0.5500 1.0500 ;
        RECT 1.5350 0.9550 2.1300 1.0550 ;
        RECT 0.3000 1.0500 0.5500 1.1500 ;
        RECT 2.0300 1.0550 2.1300 1.2500 ;
        RECT 2.0300 1.2500 2.9750 1.3500 ;
    END
    ANTENNAGATEAREA 0.3792 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.5800 3.9500 1.8200 ;
        RECT 1.6250 1.8200 3.9500 1.9200 ;
        RECT 1.6300 0.4800 3.9500 0.5800 ;
    END
    ANTENNADIFFAREA 0.87425 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 2.5300 1.6400 3.7250 1.7300 ;
      RECT 3.6350 0.7600 3.7250 1.6400 ;
      RECT 2.4300 0.6700 3.7250 0.7600 ;
      RECT 1.4750 1.2000 1.9400 1.2900 ;
      RECT 0.0650 1.3600 1.5650 1.4500 ;
      RECT 1.4750 1.2900 1.5650 1.3600 ;
      RECT 0.0650 0.7600 0.1550 1.3600 ;
      RECT 0.3550 1.4500 0.4450 1.9300 ;
      RECT 0.0650 0.6700 0.4850 0.7600 ;
      RECT 0.3150 0.4700 0.4850 0.6700 ;
      RECT 0.8900 1.6100 2.0950 1.7000 ;
      RECT 2.0050 1.5400 2.0950 1.6100 ;
      RECT 2.0050 1.4500 3.4100 1.5400 ;
      RECT 3.3200 1.0150 3.4100 1.4500 ;
      RECT 2.2300 0.9250 3.4100 1.0150 ;
      RECT 2.2300 0.7600 2.3200 0.9250 ;
      RECT 0.8500 0.6700 2.3200 0.7600 ;
      RECT 1.4100 1.7000 1.5000 1.9800 ;
      RECT 0.8900 1.7000 0.9800 1.9800 ;
      RECT 0.8500 0.4600 1.0200 0.6700 ;
  END
END XOR2_X3M_A12TH

MACRO XOR2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.5800 ;
        RECT 0.6100 0.3200 0.7100 0.6000 ;
        RECT 1.1450 0.3200 1.2450 0.5800 ;
        RECT 1.6700 0.3200 1.7600 0.5800 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.0900 1.8000 0.1900 2.0800 ;
        RECT 0.6100 1.8000 0.7100 2.0800 ;
        RECT 1.1450 1.8000 1.2450 2.0800 ;
        RECT 1.6650 1.8000 1.7650 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 1.5500 1.1500 ;
    END
    ANTENNAGATEAREA 0.3744 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5750 0.8500 2.1350 0.9500 ;
        RECT 2.0350 0.9500 2.1350 0.9550 ;
        RECT 0.5750 0.9500 0.6750 1.0450 ;
        RECT 2.0350 0.9550 2.8950 1.0550 ;
        RECT 0.2800 1.0450 0.6750 1.1450 ;
        RECT 2.7950 1.0550 2.8950 1.2500 ;
        RECT 2.7950 1.2500 4.0200 1.3500 ;
    END
    ANTENNAGATEAREA 0.4992 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 0.5800 5.5500 1.8200 ;
        RECT 1.8750 1.8200 5.5500 1.9200 ;
        RECT 1.8900 0.4800 5.5500 0.5800 ;
        RECT 2.9800 1.6300 3.1500 1.8200 ;
    END
    ANTENNADIFFAREA 1.29675 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0650 1.3600 2.0500 1.4500 ;
      RECT 1.9600 1.2900 2.0500 1.3600 ;
      RECT 1.9600 1.2000 2.6750 1.2900 ;
      RECT 0.0650 0.7600 0.1550 1.3600 ;
      RECT 0.3550 1.4500 0.4450 1.7700 ;
      RECT 0.0650 0.6700 0.4850 0.7600 ;
      RECT 0.3150 0.4700 0.4850 0.6700 ;
      RECT 2.7700 1.4450 4.6800 1.5350 ;
      RECT 4.5900 1.1200 4.6800 1.4450 ;
      RECT 4.5900 1.0300 5.0500 1.1200 ;
      RECT 4.5900 1.0150 4.6800 1.0300 ;
      RECT 2.9950 0.9250 4.6800 1.0150 ;
      RECT 2.9950 0.7600 3.0850 0.9250 ;
      RECT 0.8500 0.6700 3.0850 0.7600 ;
      RECT 0.8900 1.5700 2.8600 1.6600 ;
      RECT 2.7700 1.5350 2.8600 1.5700 ;
      RECT 0.8900 1.6600 0.9800 1.9700 ;
      RECT 0.8500 0.4700 1.0200 0.6700 ;
      RECT 1.4100 1.6600 1.5000 1.9600 ;
      RECT 1.3700 0.4700 1.5400 0.6700 ;
      RECT 3.3000 1.6400 5.2600 1.7300 ;
      RECT 5.1700 0.7600 5.2600 1.6400 ;
      RECT 3.1950 0.6700 5.2600 0.7600 ;
  END
END XOR2_X4M_A12TH

MACRO XOR3_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6750 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.7500 1.5500 ;
        RECT 0.6500 1.5500 0.7500 1.8200 ;
        RECT 0.2500 1.1400 0.3500 1.4500 ;
        RECT 0.6500 1.8200 1.5100 1.9200 ;
        RECT 0.2500 1.0400 0.9600 1.1400 ;
        RECT 1.3400 1.9200 1.5100 1.9850 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6300 0.5750 3.7500 1.9700 ;
    END
    ANTENNADIFFAREA 0.134475 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0350 0.8600 2.1500 1.8200 ;
        RECT 2.0350 1.8200 2.9900 1.9200 ;
        RECT 2.8200 1.9200 2.9900 1.9800 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.2500 1.0000 1.3500 ;
    END
    ANTENNAGATEAREA 0.0453 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 3.3250 1.8900 3.4950 2.0800 ;
        RECT 0.3900 1.7600 0.5000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8750 0.4800 2.5300 0.5700 ;
      RECT 2.4400 0.5700 2.5300 0.6800 ;
      RECT 2.4400 0.6800 2.8350 0.7700 ;
      RECT 2.7450 0.7700 2.8350 1.0500 ;
      RECT 2.7450 1.0500 3.1800 1.1400 ;
      RECT 2.7450 1.1400 2.8350 1.4300 ;
      RECT 2.4900 1.4300 2.8350 1.5200 ;
      RECT 2.4900 1.5200 2.5800 1.6550 ;
      RECT 1.1350 1.6400 1.8750 1.7300 ;
      RECT 1.7850 0.5700 1.8750 1.6400 ;
      RECT 2.9850 1.4600 3.3600 1.5500 ;
      RECT 3.2700 0.7700 3.3600 1.4600 ;
      RECT 2.9450 0.6800 3.3600 0.7700 ;
      RECT 2.7050 1.6400 3.5400 1.7300 ;
      RECT 3.4500 0.5900 3.5400 1.6400 ;
      RECT 2.6550 0.5000 3.5400 0.5900 ;
      RECT 0.0500 0.8400 1.1800 0.9300 ;
      RECT 1.0900 0.9300 1.1800 1.0750 ;
      RECT 0.0500 1.6600 0.2450 1.7500 ;
      RECT 0.0500 0.9300 0.1400 1.6600 ;
      RECT 0.0500 0.5550 0.1700 0.8400 ;
      RECT 0.9100 1.5450 1.0000 1.6800 ;
      RECT 0.9100 1.4550 1.4100 1.5450 ;
      RECT 1.3200 0.7500 1.4100 1.4550 ;
      RECT 0.6200 0.6600 1.4100 0.7500 ;
      RECT 1.5000 0.7500 1.5900 1.5300 ;
      RECT 1.5000 0.6600 1.6700 0.7500 ;
      RECT 2.2400 1.3100 2.3300 1.5650 ;
      RECT 2.2400 1.2200 2.5950 1.3100 ;
      RECT 2.5050 0.9700 2.5950 1.2200 ;
      RECT 2.2400 0.8800 2.5950 0.9700 ;
      RECT 2.2400 0.7500 2.3300 0.8800 ;
      RECT 2.1150 0.6600 2.3300 0.7500 ;
  END
END XOR3_X0P5M_A12TH

MACRO SDFFRPQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 1.0000 0.3200 1.1000 0.7350 ;
        RECT 5.6750 0.3200 5.8450 0.8400 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.3950 1.4600 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END SE

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.2850 1.7100 ;
        RECT 5.1850 0.7700 5.2850 1.4100 ;
        RECT 5.1150 0.6800 5.2850 0.7700 ;
    END
    ANTENNADIFFAREA 0.143075 ;
  END QN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.1500 2.5500 1.3900 ;
        RECT 2.4500 1.0500 2.7200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0537 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.9900 1.7300 1.1600 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3750 1.0700 1.5550 1.4400 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0250 0.9500 1.4450 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.0050 5.9250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.0600 1.8300 0.7450 1.9200 ;
      RECT 0.0600 0.5600 0.5750 0.6500 ;
      RECT 0.4850 0.5000 0.5750 0.5600 ;
      RECT 0.4850 0.4100 0.7900 0.5000 ;
      RECT 0.0600 0.6500 0.1500 1.8300 ;
      RECT 1.4700 1.6400 1.5800 1.7800 ;
      RECT 0.4550 1.5400 1.5800 1.6400 ;
      RECT 0.4100 0.8350 1.5900 0.9250 ;
      RECT 1.4900 0.5650 1.5900 0.8350 ;
      RECT 1.1050 0.9250 1.1950 1.5400 ;
      RECT 1.9050 0.8500 2.9500 0.9400 ;
      RECT 2.8600 0.9400 2.9500 1.3800 ;
      RECT 1.7450 1.5750 1.9950 1.6650 ;
      RECT 1.9050 0.9400 1.9950 1.5750 ;
      RECT 1.9050 0.6700 1.9950 0.8500 ;
      RECT 2.1750 1.5700 3.1900 1.6600 ;
      RECT 3.1000 0.7500 3.1900 1.5700 ;
      RECT 2.6950 0.6600 3.1900 0.7500 ;
      RECT 2.1750 1.2400 2.2650 1.5700 ;
      RECT 4.4550 1.1900 4.6500 1.3000 ;
      RECT 4.4550 1.0600 4.5450 1.1900 ;
      RECT 4.0350 0.9900 4.5450 1.0600 ;
      RECT 3.3350 0.9700 4.5450 0.9900 ;
      RECT 3.3350 0.9900 3.4250 1.6950 ;
      RECT 3.3350 0.9000 4.1250 0.9700 ;
      RECT 3.8550 1.5350 4.8850 1.6250 ;
      RECT 3.8550 1.2350 3.9450 1.5350 ;
      RECT 4.7950 0.7800 4.8850 1.5350 ;
      RECT 4.4250 0.6700 4.8850 0.7800 ;
      RECT 1.7050 0.4800 5.5200 0.5700 ;
      RECT 5.4300 0.5700 5.5200 1.7100 ;
      RECT 1.7050 0.5700 1.7950 1.4750 ;
      RECT 1.8750 1.8300 6.1200 1.9200 ;
      RECT 6.0300 0.7000 6.1200 1.8300 ;
      RECT 3.5850 1.1100 3.6750 1.8300 ;
  END
END SDFFRPQN_X0P5M_A12TH

MACRO SDFFRPQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0600 0.3200 0.2000 0.4650 ;
        RECT 1.0050 0.3200 1.1050 0.5100 ;
        RECT 5.7150 0.3200 5.8150 0.8750 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.2800 1.6500 ;
        RECT 5.1800 0.6800 5.2800 1.4100 ;
    END
    ANTENNADIFFAREA 0.248 ;
  END QN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0500 0.3900 1.4600 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6450 1.0050 2.9050 1.1950 ;
    END
    ANTENNAGATEAREA 0.0864 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.9950 1.9650 1.1250 2.0800 ;
        RECT 0.1050 1.8650 0.2150 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0800 1.4500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.0550 0.9500 1.5100 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6450 1.0050 5.8950 1.2050 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3150 1.8800 0.7300 1.9700 ;
      RECT 0.3150 1.7200 0.4050 1.8800 ;
      RECT 0.0600 1.6300 0.4050 1.7200 ;
      RECT 0.0600 0.6000 0.4900 0.6900 ;
      RECT 0.4000 0.5100 0.4900 0.6000 ;
      RECT 0.4000 0.4200 0.7700 0.5100 ;
      RECT 0.0600 0.6900 0.1500 1.6300 ;
      RECT 1.0600 1.7450 1.6100 1.7900 ;
      RECT 0.4950 1.7000 1.6100 1.7450 ;
      RECT 0.4400 0.8550 1.5500 0.9450 ;
      RECT 1.4600 0.6300 1.5500 0.8550 ;
      RECT 0.4950 1.6550 1.1500 1.7000 ;
      RECT 1.0600 0.9450 1.1500 1.6550 ;
      RECT 0.4950 1.5450 0.5850 1.6550 ;
      RECT 0.4400 0.8350 0.6250 0.8550 ;
      RECT 1.7000 1.6150 1.9300 1.7050 ;
      RECT 1.8400 1.0800 1.9300 1.6150 ;
      RECT 1.8400 0.9900 2.5350 1.0800 ;
      RECT 2.4250 1.0800 2.5350 1.1650 ;
      RECT 1.8400 0.6800 1.9300 0.9900 ;
      RECT 2.0900 1.6150 2.9900 1.7050 ;
      RECT 2.9000 1.4550 2.9900 1.6150 ;
      RECT 2.9000 1.3650 3.1100 1.4550 ;
      RECT 3.0200 0.9850 3.1100 1.3650 ;
      RECT 3.0200 0.8950 3.6550 0.9850 ;
      RECT 3.0200 0.8250 3.1100 0.8950 ;
      RECT 2.5850 0.7350 3.1100 0.8250 ;
      RECT 2.0900 1.2550 2.1800 1.6150 ;
      RECT 3.1200 1.5750 3.8550 1.6650 ;
      RECT 3.7650 0.8000 3.8550 1.5750 ;
      RECT 3.2250 0.7100 4.5850 0.8000 ;
      RECT 4.4950 0.8000 4.5850 1.2400 ;
      RECT 4.2100 1.5450 4.8550 1.6350 ;
      RECT 4.2100 1.0750 4.3000 1.5450 ;
      RECT 4.7650 0.8150 4.8550 1.5450 ;
      RECT 4.6850 0.7250 4.8550 0.8150 ;
      RECT 1.6400 0.4850 5.5250 0.5750 ;
      RECT 5.4350 0.5750 5.5250 1.5000 ;
      RECT 1.6400 0.5750 1.7300 1.4900 ;
      RECT 1.8400 1.8950 6.1150 1.9200 ;
      RECT 2.0650 1.8300 6.1150 1.8950 ;
      RECT 6.0250 0.6900 6.1150 1.8300 ;
      RECT 3.9750 0.9200 4.0650 1.8300 ;
      RECT 1.8400 1.9200 2.1550 1.9850 ;
  END
END SDFFRPQN_X1M_A12TH

MACRO SDFFRPQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0750 0.3200 0.2150 0.4650 ;
        RECT 1.0450 0.3200 1.1450 0.6900 ;
        RECT 6.0700 0.3200 6.1700 0.8700 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4200 1.4800 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6950 1.0050 2.9850 1.1950 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.0850 1.8750 0.2050 2.0800 ;
        RECT 1.0200 1.8400 1.1400 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3800 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.087 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2250 0.7350 5.3500 1.7000 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0400 0.9600 1.4600 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0000 1.0100 6.2450 1.2000 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8800 0.7550 1.9700 ;
      RECT 0.3400 1.7650 0.4300 1.8800 ;
      RECT 0.0600 1.6750 0.4300 1.7650 ;
      RECT 0.0600 0.6000 0.5150 0.6900 ;
      RECT 0.4250 0.5000 0.5150 0.6000 ;
      RECT 0.4250 0.4100 0.7950 0.5000 ;
      RECT 0.0600 0.6900 0.1500 1.6750 ;
      RECT 0.5200 1.6250 1.6300 1.7150 ;
      RECT 0.4800 0.8450 1.6050 0.9350 ;
      RECT 1.5150 0.5250 1.6050 0.8450 ;
      RECT 1.1300 0.9350 1.2200 1.6250 ;
      RECT 0.5200 1.5450 0.6100 1.6250 ;
      RECT 1.7200 1.5850 1.9750 1.6750 ;
      RECT 1.8850 1.1900 1.9750 1.5850 ;
      RECT 1.8850 1.1000 2.5950 1.1900 ;
      RECT 2.4850 0.9750 2.5950 1.1000 ;
      RECT 1.8850 0.7000 1.9750 1.1000 ;
      RECT 2.8700 1.4250 2.9600 1.7250 ;
      RECT 2.0750 1.3350 3.6500 1.4250 ;
      RECT 3.5600 0.9200 3.6500 1.3350 ;
      RECT 3.1150 0.8300 3.2050 1.3350 ;
      RECT 2.6350 0.7400 3.2050 0.8300 ;
      RECT 3.1050 1.5950 3.9100 1.6850 ;
      RECT 3.8200 0.7900 3.9100 1.5950 ;
      RECT 3.3300 0.7000 4.6050 0.7900 ;
      RECT 3.3300 0.7900 3.4200 0.8700 ;
      RECT 4.5150 0.7900 4.6050 1.2750 ;
      RECT 4.2450 1.5550 4.8750 1.6450 ;
      RECT 4.2450 1.1100 4.3350 1.5550 ;
      RECT 4.7850 0.8150 4.8750 1.5550 ;
      RECT 4.7050 0.7250 4.8750 0.8150 ;
      RECT 1.6950 0.4900 5.8600 0.5800 ;
      RECT 5.7600 0.5800 5.8600 1.6700 ;
      RECT 1.6600 1.2850 1.7850 1.4550 ;
      RECT 1.6950 0.5800 1.7850 1.2850 ;
      RECT 1.9900 0.4100 2.0800 0.4900 ;
      RECT 1.8950 1.8300 6.4800 1.9200 ;
      RECT 6.3900 0.6850 6.4800 1.8300 ;
      RECT 3.0500 1.9200 3.2200 1.9450 ;
      RECT 4.0100 0.9300 4.1000 1.8300 ;
      RECT 1.8950 1.9200 2.0650 1.9850 ;
  END
END SDFFRPQN_X2M_A12TH

MACRO SDFFRPQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.0800 0.3200 0.2100 0.4650 ;
        RECT 1.0350 0.3200 1.1550 0.6500 ;
        RECT 5.4450 0.3200 5.5450 0.6800 ;
        RECT 5.9450 0.3200 6.1150 0.5150 ;
        RECT 6.5000 0.3200 6.6000 0.6250 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0850 0.4200 1.4550 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7200 1.0050 2.9750 1.1950 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 4.4300 2.0400 4.6000 2.0800 ;
        RECT 5.9850 2.0350 6.0750 2.0800 ;
        RECT 6.4650 1.8850 6.6350 2.0800 ;
        RECT 1.0350 1.8400 1.1550 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0500 1.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2450 1.6500 6.8550 1.7500 ;
        RECT 6.7650 1.7500 6.8550 1.9150 ;
        RECT 6.2450 0.5400 6.3350 1.6500 ;
        RECT 6.7650 0.5400 6.8550 1.6500 ;
    END
    ANTENNADIFFAREA 0.58175 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0400 0.9600 1.4500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6300 1.0100 5.8500 1.2050 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3350 1.8800 0.7500 1.9700 ;
      RECT 0.3350 1.7600 0.4250 1.8800 ;
      RECT 0.0600 1.6700 0.4250 1.7600 ;
      RECT 0.0600 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5050 0.5100 0.6000 ;
      RECT 0.4200 0.4150 0.7900 0.5050 ;
      RECT 0.0600 0.6900 0.1500 1.6700 ;
      RECT 1.4750 1.7150 1.6450 1.9700 ;
      RECT 0.5150 1.6250 1.6450 1.7150 ;
      RECT 0.4750 0.8550 1.6050 0.9450 ;
      RECT 1.5150 0.6700 1.6050 0.8550 ;
      RECT 1.1350 0.9450 1.2250 1.6250 ;
      RECT 0.5150 1.5450 0.6050 1.6250 ;
      RECT 0.4750 0.8150 0.6450 0.8550 ;
      RECT 1.7350 1.5800 1.9750 1.6700 ;
      RECT 1.8850 1.1650 1.9750 1.5800 ;
      RECT 1.8850 1.0750 2.5500 1.1650 ;
      RECT 2.4500 0.9750 2.5500 1.0750 ;
      RECT 1.8850 0.7000 1.9750 1.0750 ;
      RECT 2.1500 1.4950 3.0300 1.5850 ;
      RECT 2.9400 1.4550 3.0300 1.4950 ;
      RECT 2.9400 1.3650 3.7350 1.4550 ;
      RECT 3.6450 0.9200 3.7350 1.3650 ;
      RECT 3.1250 0.8300 3.2150 1.3650 ;
      RECT 2.6900 0.7400 3.2150 0.8300 ;
      RECT 2.1500 1.2650 2.2400 1.4950 ;
      RECT 3.1700 1.5950 3.9950 1.6850 ;
      RECT 3.9050 0.7900 3.9950 1.5950 ;
      RECT 3.3650 0.7000 4.7450 0.7900 ;
      RECT 3.3650 0.7900 3.4700 0.8750 ;
      RECT 4.6550 0.7900 4.7450 1.1950 ;
      RECT 4.3650 1.4100 4.9800 1.5000 ;
      RECT 4.3650 0.9100 4.4550 1.4100 ;
      RECT 4.8900 0.6750 4.9800 1.4100 ;
      RECT 1.6950 0.4900 5.2400 0.5800 ;
      RECT 5.1500 0.5800 5.2400 1.4700 ;
      RECT 1.6600 1.3000 1.7850 1.4700 ;
      RECT 1.6950 0.5800 1.7850 1.3000 ;
      RECT 2.0150 0.4100 2.1050 0.4900 ;
      RECT 5.4000 1.5000 5.8950 1.5900 ;
      RECT 5.4000 0.7900 5.8550 0.8800 ;
      RECT 5.7650 0.6750 5.8550 0.7900 ;
      RECT 4.1300 1.6200 5.4900 1.7100 ;
      RECT 5.4000 1.5900 5.4900 1.6200 ;
      RECT 5.4000 0.8800 5.4900 1.5000 ;
      RECT 1.8750 1.8800 4.2200 1.9200 ;
      RECT 2.1100 1.8300 4.2200 1.8800 ;
      RECT 4.1300 1.7100 4.2200 1.8300 ;
      RECT 4.1300 0.9300 4.2200 1.6200 ;
      RECT 1.8750 1.9200 2.2000 1.9700 ;
      RECT 4.6950 1.8300 6.1400 1.9200 ;
      RECT 6.0500 1.0100 6.1400 1.8300 ;
  END
END SDFFRPQN_X3M_A12TH

MACRO SDFFRPQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6900 ;
        RECT 1.0300 0.3200 1.1300 0.7300 ;
        RECT 5.7100 0.3200 5.8100 0.8850 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1800 1.5100 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.2800 1.7100 ;
        RECT 5.1800 0.6700 5.2800 1.4100 ;
    END
    ANTENNADIFFAREA 0.1322 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.1550 2.5500 1.3900 ;
        RECT 2.4500 1.0550 2.7450 1.1550 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.0900 1.8150 0.1900 2.0800 ;
        RECT 1.0250 1.7900 1.1250 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0700 1.5500 1.4400 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0500 0.9550 1.4700 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.0050 5.9250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3300 1.8300 0.7450 1.9200 ;
      RECT 0.3300 1.7700 0.4200 1.8300 ;
      RECT 0.2800 1.6800 0.4200 1.7700 ;
      RECT 0.2800 0.7250 0.3700 1.6800 ;
      RECT 0.2800 0.6350 0.5050 0.7250 ;
      RECT 0.4150 0.5200 0.5050 0.6350 ;
      RECT 0.4150 0.4300 0.8050 0.5200 ;
      RECT 0.5100 1.6000 1.6450 1.7000 ;
      RECT 0.4700 0.8350 1.5900 0.9250 ;
      RECT 1.4900 0.7450 1.5900 0.8350 ;
      RECT 1.0550 0.9250 1.1450 1.6000 ;
      RECT 0.5100 1.5200 0.6000 1.6000 ;
      RECT 1.9300 0.8500 2.9750 0.9400 ;
      RECT 2.8850 0.9400 2.9750 1.2400 ;
      RECT 2.8800 1.2400 2.9750 1.4100 ;
      RECT 1.7700 1.5750 2.0200 1.6650 ;
      RECT 1.9300 0.9400 2.0200 1.5750 ;
      RECT 1.9300 0.6700 2.0200 0.8500 ;
      RECT 2.1850 1.5700 3.1900 1.6600 ;
      RECT 3.1000 0.7500 3.1900 1.5700 ;
      RECT 2.7150 0.6600 3.1900 0.7500 ;
      RECT 2.1850 1.2600 2.2750 1.5700 ;
      RECT 4.3800 1.1900 4.5850 1.3000 ;
      RECT 4.3800 0.7850 4.4700 1.1900 ;
      RECT 3.3350 0.6950 4.4700 0.7850 ;
      RECT 3.3350 0.7850 3.4250 1.6950 ;
      RECT 4.7950 1.0550 5.0650 1.1450 ;
      RECT 3.8700 1.5500 4.8850 1.6400 ;
      RECT 4.7950 1.1450 4.8850 1.5500 ;
      RECT 3.8700 1.0100 3.9600 1.5500 ;
      RECT 4.7950 0.9400 4.8850 1.0550 ;
      RECT 4.5650 0.8300 4.8850 0.9400 ;
      RECT 4.5650 0.6700 4.6750 0.8300 ;
      RECT 1.7100 0.4800 5.5200 0.5700 ;
      RECT 5.4300 0.5700 5.5200 1.7100 ;
      RECT 1.7100 1.2850 1.8150 1.4550 ;
      RECT 1.7100 0.5700 1.8000 1.2850 ;
      RECT 1.8950 1.8300 6.1200 1.9200 ;
      RECT 6.0300 0.7000 6.1200 1.8300 ;
      RECT 3.6150 1.0950 3.7050 1.8300 ;
  END
END SDFFRPQ_X0P5M_A12TH

MACRO SDFFRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4650 ;
        RECT 1.0550 0.3200 1.1550 0.6750 ;
        RECT 5.9050 0.3200 6.0050 0.8450 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1700 1.4600 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 1.4100 5.4400 1.6500 ;
        RECT 5.3400 0.7050 5.4400 1.4100 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.0500 3.0600 1.1500 ;
    END
    ANTENNAGATEAREA 0.093 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 2.3550 2.0650 2.5250 2.0800 ;
        RECT 5.9100 1.9650 6.0000 2.0800 ;
        RECT 4.3700 1.9400 4.5400 2.0800 ;
        RECT 1.0150 1.9350 1.1850 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9500 1.4750 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 1.0000 6.0900 1.1900 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3300 1.8800 0.7400 1.9700 ;
      RECT 0.3300 1.8600 0.4200 1.8800 ;
      RECT 0.2750 1.7700 0.4200 1.8600 ;
      RECT 0.2750 0.6900 0.3650 1.7700 ;
      RECT 0.2750 0.6000 0.5000 0.6900 ;
      RECT 0.4100 0.5200 0.5000 0.6000 ;
      RECT 0.4100 0.4300 0.7800 0.5200 ;
      RECT 0.5050 1.6250 1.6500 1.7150 ;
      RECT 0.5050 0.8000 1.6100 0.8900 ;
      RECT 1.5200 0.4800 1.6100 0.8000 ;
      RECT 1.0550 0.8900 1.1450 1.6250 ;
      RECT 0.5050 1.5450 0.5950 1.6250 ;
      RECT 0.5050 0.8900 0.5950 1.0050 ;
      RECT 1.7400 1.6150 1.9800 1.7050 ;
      RECT 1.8900 1.1900 1.9800 1.6150 ;
      RECT 1.8900 1.1000 2.5500 1.1900 ;
      RECT 2.4500 0.9700 2.5500 1.1000 ;
      RECT 1.8900 0.7100 1.9800 1.1000 ;
      RECT 2.1300 1.5950 3.0250 1.6850 ;
      RECT 2.9350 1.4550 3.0250 1.5950 ;
      RECT 2.9350 1.3650 3.2600 1.4550 ;
      RECT 3.1700 1.1000 3.2600 1.3650 ;
      RECT 3.1700 1.0100 3.6700 1.1000 ;
      RECT 3.5800 0.9850 3.6700 1.0100 ;
      RECT 3.1700 0.8500 3.2600 1.0100 ;
      RECT 3.5800 0.8950 3.7900 0.9850 ;
      RECT 2.6900 0.7600 3.2600 0.8500 ;
      RECT 2.1300 1.3000 2.2200 1.5950 ;
      RECT 3.1350 1.5950 3.9900 1.6850 ;
      RECT 3.9000 0.8000 3.9900 1.5950 ;
      RECT 3.3600 0.7100 4.7300 0.8000 ;
      RECT 3.3600 0.8000 3.4500 0.9000 ;
      RECT 4.6400 0.8000 4.7300 1.0800 ;
      RECT 4.6400 1.0800 4.8150 1.2850 ;
      RECT 4.3750 1.5500 5.0200 1.6400 ;
      RECT 4.9300 1.1700 5.0200 1.5500 ;
      RECT 4.3750 0.9200 4.4650 1.5500 ;
      RECT 4.9300 1.0800 5.1400 1.1700 ;
      RECT 4.9300 0.7700 5.0200 1.0800 ;
      RECT 4.8400 0.6800 5.0200 0.7700 ;
      RECT 1.7000 0.4850 5.7150 0.5750 ;
      RECT 5.6250 0.5750 5.7150 1.4800 ;
      RECT 1.6550 1.3250 1.7900 1.4950 ;
      RECT 1.7000 0.5750 1.7900 1.3250 ;
      RECT 2.1050 1.8300 6.3050 1.8400 ;
      RECT 4.1300 1.7500 6.3050 1.8300 ;
      RECT 6.2150 0.6400 6.3050 1.7500 ;
      RECT 1.8250 1.8950 4.2200 1.9200 ;
      RECT 2.1050 1.8400 4.2200 1.8950 ;
      RECT 4.1300 0.9300 4.2200 1.7500 ;
      RECT 1.8250 1.9200 2.1950 1.9850 ;
  END
END SDFFRPQ_X1M_A12TH

MACRO SDFFRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.6900 ;
        RECT 1.0600 0.3200 1.2000 0.6900 ;
        RECT 6.1050 0.3200 6.2050 0.9050 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0700 0.1700 1.6100 ;
    END
    ANTENNAGATEAREA 0.0684 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9500 1.4300 ;
    END
    ANTENNAGATEAREA 0.102 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.0900 1.8650 0.2000 2.0800 ;
        RECT 1.0650 1.8300 1.1850 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4300 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2450 1.4100 5.3950 1.6950 ;
        RECT 5.2950 0.7050 5.3950 1.4100 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0400 0.9900 1.4500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0400 1.0100 6.3150 1.1900 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8800 0.7550 1.9700 ;
      RECT 0.3400 1.8300 0.4300 1.8800 ;
      RECT 0.2900 1.7400 0.4300 1.8300 ;
      RECT 0.2900 0.6700 0.3800 1.7400 ;
      RECT 0.2900 0.5800 0.5150 0.6700 ;
      RECT 0.4250 0.5200 0.5150 0.5800 ;
      RECT 0.4250 0.4300 0.8150 0.5200 ;
      RECT 0.5200 1.6400 1.6700 1.7300 ;
      RECT 0.4950 0.8150 1.6300 0.9050 ;
      RECT 1.5400 0.4950 1.6300 0.8150 ;
      RECT 1.0900 0.9050 1.1800 1.6400 ;
      RECT 0.5200 1.5450 0.6100 1.6400 ;
      RECT 1.7700 1.5950 2.0150 1.6850 ;
      RECT 1.9250 1.1500 2.0150 1.5950 ;
      RECT 1.9250 1.0600 2.6900 1.1500 ;
      RECT 2.5800 0.9600 2.6900 1.0600 ;
      RECT 1.9250 0.6800 2.0150 1.0600 ;
      RECT 2.2500 1.5950 3.2050 1.6850 ;
      RECT 3.1150 1.1100 3.2050 1.5950 ;
      RECT 3.1150 1.0200 3.7150 1.1100 ;
      RECT 3.6150 0.9000 3.7150 1.0200 ;
      RECT 3.1150 0.8300 3.2050 1.0200 ;
      RECT 2.6950 0.7400 3.2050 0.8300 ;
      RECT 2.2500 1.2700 2.3400 1.5950 ;
      RECT 3.3250 1.5950 3.9700 1.6850 ;
      RECT 3.8800 0.7850 3.9700 1.5950 ;
      RECT 3.3700 0.6950 4.6400 0.7850 ;
      RECT 3.3700 0.7850 3.4600 0.8850 ;
      RECT 4.5500 0.7850 4.6400 0.9250 ;
      RECT 4.5500 0.9250 4.6850 1.0150 ;
      RECT 4.5950 1.0150 4.6850 1.3500 ;
      RECT 4.3500 1.5650 4.9550 1.6550 ;
      RECT 4.8650 1.1800 4.9550 1.5650 ;
      RECT 4.3500 1.0850 4.4400 1.5650 ;
      RECT 4.8650 1.0700 5.1500 1.1800 ;
      RECT 4.8650 0.8300 4.9550 1.0700 ;
      RECT 4.7550 0.7200 4.9550 0.8300 ;
      RECT 1.7250 0.4900 5.8700 0.5800 ;
      RECT 5.7800 0.5800 5.8700 1.6900 ;
      RECT 1.7250 0.5800 1.8150 1.4850 ;
      RECT 2.0500 0.4100 2.1400 0.4900 ;
      RECT 1.9500 1.8300 6.1450 1.9200 ;
      RECT 6.0550 1.5350 6.1450 1.8300 ;
      RECT 6.0550 1.4450 6.5450 1.5350 ;
      RECT 6.4550 0.8500 6.5450 1.4450 ;
      RECT 6.3550 0.7600 6.5450 0.8500 ;
      RECT 4.1100 0.9100 4.2000 1.8300 ;
  END
END SDFFRPQ_X2M_A12TH

MACRO SDFFRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7200 ;
        RECT 1.0350 0.3200 1.1550 0.6750 ;
        RECT 6.3550 0.3200 6.4450 0.6100 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0850 0.1700 1.5450 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7100 1.0050 2.9700 1.1950 ;
    END
    ANTENNAGATEAREA 0.0981 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 0.0950 1.8650 0.1950 2.0800 ;
        RECT 1.0350 1.8400 1.1550 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.0850 1.5500 1.5050 ;
    END
    ANTENNAGATEAREA 0.0882 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0950 1.2500 6.7100 1.3500 ;
        RECT 6.0950 1.3500 6.1850 1.7000 ;
        RECT 6.6100 1.3500 6.7100 1.7000 ;
        RECT 6.6100 0.9500 6.7100 1.2500 ;
        RECT 6.0900 0.8500 6.7100 0.9500 ;
        RECT 6.0900 0.4850 6.1900 0.8500 ;
        RECT 6.6100 0.4850 6.7100 0.8500 ;
    END
    ANTENNADIFFAREA 0.595725 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0400 0.9700 1.4500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4400 1.0100 5.7000 1.1900 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3350 1.8800 0.7500 1.9700 ;
      RECT 0.3350 1.8200 0.4250 1.8800 ;
      RECT 0.2850 1.7300 0.4250 1.8200 ;
      RECT 0.2850 0.7000 0.3750 1.7300 ;
      RECT 0.2850 0.6100 0.5100 0.7000 ;
      RECT 0.4200 0.5300 0.5100 0.6100 ;
      RECT 0.4200 0.4400 0.8200 0.5300 ;
      RECT 1.4750 1.7300 1.6450 1.9700 ;
      RECT 0.5150 1.6400 1.6450 1.7300 ;
      RECT 0.4750 0.8550 1.6050 0.9450 ;
      RECT 1.5150 0.5350 1.6050 0.8550 ;
      RECT 1.0600 0.9450 1.1500 1.6400 ;
      RECT 0.5150 1.5450 0.6050 1.6400 ;
      RECT 1.7350 1.6150 1.9650 1.7050 ;
      RECT 1.8750 1.1900 1.9650 1.6150 ;
      RECT 1.8750 1.1000 2.5600 1.1900 ;
      RECT 2.4400 0.9900 2.5600 1.1000 ;
      RECT 1.8750 0.7000 1.9650 1.1000 ;
      RECT 2.1100 1.5950 3.1700 1.6850 ;
      RECT 3.0800 1.0500 3.1700 1.5950 ;
      RECT 3.0800 0.9600 3.7000 1.0500 ;
      RECT 3.0800 0.8300 3.1700 0.9600 ;
      RECT 2.6150 0.7400 3.1700 0.8300 ;
      RECT 2.1100 1.2950 2.2000 1.5950 ;
      RECT 3.2650 1.2800 3.3550 1.7200 ;
      RECT 3.2650 1.1900 3.8950 1.2800 ;
      RECT 3.8050 0.7900 3.8950 1.1900 ;
      RECT 3.2800 0.7000 4.3150 0.7900 ;
      RECT 3.2800 0.7900 3.4000 0.8700 ;
      RECT 4.2250 0.7900 4.3150 1.0550 ;
      RECT 4.2250 1.0550 4.7050 1.1450 ;
      RECT 1.6950 0.4900 4.5250 0.5800 ;
      RECT 4.4350 0.5800 4.5250 0.6800 ;
      RECT 4.4350 0.6800 5.0650 0.7700 ;
      RECT 4.9750 0.7700 5.0650 1.4700 ;
      RECT 1.6600 1.3000 1.7850 1.4700 ;
      RECT 1.6950 0.5800 1.7850 1.3000 ;
      RECT 1.9850 0.4100 2.0750 0.4900 ;
      RECT 5.1800 1.4600 5.7650 1.5500 ;
      RECT 5.1800 0.7300 5.7650 0.8200 ;
      RECT 1.8750 1.8800 3.7800 1.9200 ;
      RECT 3.6100 1.9200 3.7800 1.9450 ;
      RECT 2.1100 1.8300 3.7800 1.8800 ;
      RECT 3.6100 1.6800 3.7000 1.8300 ;
      RECT 3.6100 1.5900 5.2700 1.6800 ;
      RECT 5.1800 1.5500 5.2700 1.5900 ;
      RECT 4.0300 0.9400 4.1200 1.5900 ;
      RECT 5.1800 0.8200 5.2700 1.4600 ;
      RECT 1.8750 1.9200 2.2000 1.9700 ;
      RECT 5.9000 1.0500 6.3900 1.1500 ;
      RECT 3.9400 1.8150 5.9900 1.9050 ;
      RECT 5.9000 1.1500 5.9900 1.8150 ;
      RECT 5.9000 0.5700 5.9900 1.0500 ;
      RECT 4.6550 0.4800 5.9900 0.5700 ;
      RECT 3.9400 1.9050 4.0300 1.9850 ;
  END
END SDFFRPQ_X3M_A12TH

MACRO SDFFRPQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6100 ;
        RECT 1.0400 0.3200 1.1400 0.5600 ;
        RECT 1.5650 0.3200 1.6850 0.5000 ;
        RECT 5.4350 0.3200 5.6050 0.3700 ;
        RECT 5.9600 0.3200 6.1300 0.3700 ;
        RECT 7.1200 0.3200 7.2900 0.3700 ;
        RECT 7.6750 0.3200 7.7750 0.6100 ;
        RECT 8.1950 0.3200 8.2950 0.6100 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0450 0.1700 1.4400 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9600 1.2100 2.3300 1.3500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.9400 3.8400 1.1900 ;
    END
    ANTENNAGATEAREA 0.0981 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.4450 2.7200 ;
        RECT 3.2650 2.0550 3.4350 2.0800 ;
        RECT 6.5600 2.0300 6.6500 2.0800 ;
        RECT 5.4100 2.0050 5.5800 2.0800 ;
        RECT 5.9300 2.0050 6.1000 2.0800 ;
        RECT 1.5500 1.9550 1.6800 2.0800 ;
        RECT 0.1450 1.8600 0.2350 2.0800 ;
        RECT 7.6750 1.7900 7.7750 2.0800 ;
        RECT 8.1950 1.7900 8.2950 2.0800 ;
        RECT 1.0300 1.7600 1.1300 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4150 0.8500 8.1500 0.9500 ;
        RECT 8.0500 0.9500 8.1500 1.2900 ;
        RECT 7.4150 0.5000 7.5150 0.8500 ;
        RECT 7.9350 0.5000 8.0350 0.8500 ;
        RECT 7.4150 1.2900 8.1500 1.3900 ;
        RECT 7.4150 1.3900 7.5150 1.7250 ;
        RECT 7.9350 1.3900 8.0350 1.7250 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0100 0.9600 1.4200 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.7400 1.0100 6.9600 1.2150 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 4.1050 1.5950 4.3600 1.6850 ;
      RECT 4.2700 1.3250 4.3600 1.5950 ;
      RECT 4.2700 1.2350 4.9450 1.3250 ;
      RECT 4.8550 0.7900 4.9450 1.2350 ;
      RECT 4.2750 0.7000 5.3900 0.7900 ;
      RECT 5.3000 0.7900 5.3900 1.0900 ;
      RECT 5.3000 1.0900 5.9600 1.1800 ;
      RECT 6.1800 1.3250 6.3150 1.4950 ;
      RECT 6.1800 0.8750 6.2700 1.3250 ;
      RECT 6.1800 0.7950 6.3500 0.8750 ;
      RECT 5.4950 0.7050 6.3500 0.7950 ;
      RECT 5.4950 0.5700 5.5850 0.7050 ;
      RECT 2.5350 0.4800 5.5850 0.5700 ;
      RECT 4.3850 0.4500 4.5550 0.4800 ;
      RECT 2.5350 0.5700 2.6250 1.4200 ;
      RECT 2.7700 0.4400 2.9950 0.4800 ;
      RECT 6.4700 1.5050 7.0300 1.5950 ;
      RECT 6.4700 0.7500 7.0300 0.8400 ;
      RECT 2.7650 1.8800 4.7250 1.9200 ;
      RECT 2.9750 1.8300 4.7250 1.8800 ;
      RECT 4.6350 1.7050 4.7250 1.8300 ;
      RECT 4.6350 1.6150 6.5600 1.7050 ;
      RECT 6.4700 1.5950 6.5600 1.6150 ;
      RECT 5.0950 0.9000 5.1850 1.6150 ;
      RECT 6.4700 0.8400 6.5600 1.5050 ;
      RECT 2.7650 1.9200 3.0650 1.9700 ;
      RECT 7.1800 1.0800 7.7500 1.1700 ;
      RECT 4.9350 1.8150 7.2750 1.9050 ;
      RECT 7.1800 1.1700 7.2700 1.8150 ;
      RECT 7.1800 0.5800 7.2700 1.0800 ;
      RECT 5.6850 0.4900 7.2700 0.5800 ;
      RECT 4.9350 1.9050 5.1050 1.9450 ;
      RECT 0.3250 1.8800 0.7400 1.9700 ;
      RECT 0.3250 1.7150 0.4150 1.8800 ;
      RECT 0.2750 1.6250 0.4150 1.7150 ;
      RECT 0.2750 0.6900 0.3650 1.6250 ;
      RECT 0.2750 0.6000 0.5250 0.6900 ;
      RECT 0.4350 0.5100 0.5250 0.6000 ;
      RECT 0.4350 0.4200 0.7800 0.5100 ;
      RECT 1.2600 0.6000 2.2350 0.6900 ;
      RECT 1.2550 1.7650 2.2450 1.8550 ;
      RECT 0.5050 1.5700 2.5050 1.6600 ;
      RECT 0.4650 0.8100 2.4450 0.9000 ;
      RECT 2.3550 0.6750 2.4450 0.8100 ;
      RECT 1.2000 0.9000 1.2900 1.5700 ;
      RECT 0.5050 1.6600 0.5950 1.7400 ;
      RECT 2.5950 1.6150 2.8450 1.7050 ;
      RECT 2.7550 1.1200 2.8450 1.6150 ;
      RECT 2.7550 1.0300 3.5100 1.1200 ;
      RECT 3.4000 0.9100 3.5100 1.0300 ;
      RECT 2.7550 0.6600 2.8450 1.0300 ;
      RECT 3.0400 1.5950 3.9200 1.6850 ;
      RECT 3.8300 1.4550 3.9200 1.5950 ;
      RECT 3.8300 1.3650 4.1000 1.4550 ;
      RECT 4.0100 1.0500 4.1000 1.3650 ;
      RECT 4.0100 0.9600 4.7450 1.0500 ;
      RECT 4.0100 0.7800 4.1000 0.9600 ;
      RECT 3.6000 0.6900 4.1000 0.7800 ;
      RECT 3.0400 1.2300 3.1300 1.5950 ;
  END
END SDFFRPQ_X4M_A12TH

MACRO SDFFSQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 1.0000 ;
        RECT 1.1150 0.3200 1.2850 0.8000 ;
        RECT 5.6250 0.3200 5.7950 0.9200 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1950 0.2800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.0100 5.8800 1.2100 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4200 1.1350 1.5900 1.3900 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.1950 1.6500 ;
        RECT 5.0950 0.8050 5.1950 1.4100 ;
    END
    ANTENNADIFFAREA 0.13475 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.2100 3.0900 1.3900 ;
    END
    ANTENNAGATEAREA 0.0486 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.6900 1.7850 5.7900 2.0800 ;
        RECT 1.0750 1.6750 1.2450 2.0800 ;
        RECT 0.1050 1.4800 0.2050 2.0800 ;
    END
  END VDD

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9700 1.1050 1.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI
  OBS
    LAYER M1 ;
      RECT 0.3700 1.7350 0.8550 1.8250 ;
      RECT 0.3700 0.5500 0.4600 1.7350 ;
      RECT 0.3700 0.4600 0.6350 0.5500 ;
      RECT 0.5700 1.4950 1.7350 1.5850 ;
      RECT 0.6200 0.8900 1.6950 0.9800 ;
      RECT 1.6050 0.6650 1.6950 0.8900 ;
      RECT 0.6200 0.9800 0.7100 1.4950 ;
      RECT 0.6200 0.7750 0.7100 0.8900 ;
      RECT 1.8250 1.4950 2.0850 1.5850 ;
      RECT 1.9950 0.9200 2.0850 1.4950 ;
      RECT 1.9950 0.8300 2.7500 0.9200 ;
      RECT 2.6600 0.9200 2.7500 1.4000 ;
      RECT 2.2850 1.5700 3.3000 1.6700 ;
      RECT 3.2000 0.9200 3.3000 1.5700 ;
      RECT 3.0300 0.8200 3.3000 0.9200 ;
      RECT 2.2850 1.1650 2.3850 1.5700 ;
      RECT 4.4150 1.3050 4.6700 1.3950 ;
      RECT 4.4150 0.9500 4.5050 1.3050 ;
      RECT 3.8550 0.8600 4.6150 0.9500 ;
      RECT 3.8550 0.9500 3.9450 1.4000 ;
      RECT 3.4200 1.5400 4.8750 1.6300 ;
      RECT 4.7850 1.1700 4.8750 1.5400 ;
      RECT 3.4200 0.7750 3.5100 1.5400 ;
      RECT 4.6150 1.0700 5.0050 1.1700 ;
      RECT 1.8150 0.5850 5.4550 0.6750 ;
      RECT 5.3650 0.6750 5.4550 1.4700 ;
      RECT 3.6250 0.6750 3.7150 1.4400 ;
      RECT 1.7600 1.2150 1.9050 1.3850 ;
      RECT 1.8150 0.6750 1.9050 1.2150 ;
      RECT 5.3950 1.5950 6.1100 1.6950 ;
      RECT 6.0100 0.7750 6.1100 1.5950 ;
      RECT 1.9100 1.7800 5.4950 1.8800 ;
      RECT 5.3950 1.6950 5.4950 1.7800 ;
  END
END SDFFSQN_X0P5M_A12TH

MACRO SDFFSQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9300 ;
        RECT 1.0950 0.3200 1.2650 0.7200 ;
        RECT 2.5600 0.3200 2.7300 0.5550 ;
        RECT 5.6550 0.3200 5.8250 0.9250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.8100 2.0400 3.0200 2.0800 ;
        RECT 1.0950 1.8350 1.2650 2.0800 ;
        RECT 0.0850 1.6800 0.1850 2.0800 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.2200 1.6700 ;
        RECT 5.1200 0.6600 5.2200 1.4100 ;
    END
    ANTENNADIFFAREA 0.2448 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.1700 5.7500 1.4950 ;
        RECT 5.6500 1.0700 5.9050 1.1700 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1700 1.5050 ;
    END
    ANTENNAGATEAREA 0.0516 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0300 1.0600 1.1500 1.4950 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0800 1.5700 1.4700 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8450 1.1850 3.0450 1.4100 ;
    END
    ANTENNAGATEAREA 0.075 ;
  END SN
  OBS
    LAYER M1 ;
      RECT 0.3500 1.8800 0.7300 1.9700 ;
      RECT 0.3500 0.6000 0.4400 1.8800 ;
      RECT 0.3500 0.5100 0.6700 0.6000 ;
      RECT 0.5950 1.6500 1.7150 1.7400 ;
      RECT 0.5550 0.8300 1.6750 0.9200 ;
      RECT 1.5850 0.7050 1.6750 0.8300 ;
      RECT 0.5950 0.9200 0.6850 1.6500 ;
      RECT 1.8050 1.6250 2.0800 1.7150 ;
      RECT 1.9900 1.1700 2.0800 1.6250 ;
      RECT 1.9900 1.0800 2.7500 1.1700 ;
      RECT 2.6600 1.1700 2.7500 1.2900 ;
      RECT 1.9900 0.7450 2.0800 1.0800 ;
      RECT 2.2500 1.6300 3.2350 1.7300 ;
      RECT 3.1350 0.7550 3.2350 1.6300 ;
      RECT 2.2500 1.2900 2.3500 1.6300 ;
      RECT 3.3450 1.6500 4.3750 1.7400 ;
      RECT 4.2400 1.5700 4.3750 1.6500 ;
      RECT 3.3950 0.7550 3.4950 1.6500 ;
      RECT 4.2400 1.1400 4.3300 1.5700 ;
      RECT 4.2400 1.0400 4.7500 1.1400 ;
      RECT 4.4300 1.3000 4.9500 1.4000 ;
      RECT 4.8500 0.8100 4.9500 1.3000 ;
      RECT 3.8150 0.7100 4.9500 0.8100 ;
      RECT 3.8150 0.8100 3.9150 1.5400 ;
      RECT 2.8500 0.4800 5.4850 0.5700 ;
      RECT 5.3850 0.5700 5.4850 1.6550 ;
      RECT 2.3500 0.6750 2.9400 0.7650 ;
      RECT 2.8500 0.5700 2.9400 0.6750 ;
      RECT 3.5850 0.5700 3.6850 1.5400 ;
      RECT 3.2650 0.4350 3.4750 0.4800 ;
      RECT 1.6800 1.3500 1.8700 1.4400 ;
      RECT 1.7800 0.6050 1.8700 1.3500 ;
      RECT 1.7800 0.5150 2.4400 0.6050 ;
      RECT 2.3500 0.6050 2.4400 0.6750 ;
      RECT 1.9050 1.8700 6.1250 1.9200 ;
      RECT 2.1250 1.8300 6.1250 1.8700 ;
      RECT 6.0250 0.7450 6.1250 1.8300 ;
      RECT 3.2450 1.9200 3.4750 1.9850 ;
      RECT 1.9050 1.9200 2.2150 1.9600 ;
  END
END SDFFSQN_X1M_A12TH

MACRO SDFFSQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9200 ;
        RECT 5.7150 0.3200 5.8150 0.8900 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9900 1.2800 5.1550 1.6500 ;
        RECT 5.0550 0.7900 5.1550 1.2800 ;
        RECT 4.9250 0.6900 5.1550 0.7900 ;
    END
    ANTENNADIFFAREA 0.306 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9750 2.9500 1.3950 ;
    END
    ANTENNAGATEAREA 0.1014 ;
  END SN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8200 1.0100 5.9500 1.3350 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.7400 2.0750 5.8300 2.0800 ;
        RECT 2.7300 2.0400 2.9000 2.0800 ;
        RECT 1.0650 1.8200 1.1650 2.0800 ;
        RECT 0.0750 1.6800 0.1750 2.0800 ;
    END
  END VDD

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2900 0.9500 1.4900 ;
        RECT 0.8500 1.1200 1.0350 1.2900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4300 1.0200 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8300 0.8050 1.9200 ;
      RECT 0.3400 0.5500 0.4300 1.8300 ;
      RECT 0.3400 0.4600 0.6150 0.5500 ;
      RECT 1.5250 1.6800 1.6250 1.9800 ;
      RECT 0.5700 1.5900 1.6250 1.6800 ;
      RECT 0.5700 0.7100 1.6400 0.8000 ;
      RECT 1.5500 0.4300 1.6400 0.7100 ;
      RECT 0.5700 0.8000 0.6600 1.5900 ;
      RECT 1.7300 1.5400 2.0350 1.6400 ;
      RECT 1.9350 0.8450 2.0350 1.5400 ;
      RECT 1.9350 0.7450 2.7100 0.8450 ;
      RECT 2.6100 0.8450 2.7100 1.2900 ;
      RECT 2.2150 1.6300 3.1400 1.7300 ;
      RECT 3.0400 0.8100 3.1400 1.6300 ;
      RECT 2.9050 0.7100 3.1400 0.8100 ;
      RECT 2.2150 1.2400 2.3150 1.6300 ;
      RECT 3.2400 1.6500 4.2350 1.7400 ;
      RECT 3.2400 1.5950 3.4350 1.6500 ;
      RECT 4.1450 1.1400 4.2350 1.6500 ;
      RECT 3.2400 0.7050 3.3300 1.5950 ;
      RECT 4.1450 1.0500 4.5500 1.1400 ;
      RECT 4.3350 1.3050 4.7900 1.3950 ;
      RECT 4.7000 0.8050 4.7900 1.3050 ;
      RECT 3.6900 0.7150 4.7900 0.8050 ;
      RECT 3.6900 0.8050 3.7800 1.5200 ;
      RECT 1.7300 0.4800 5.5500 0.5700 ;
      RECT 5.4500 0.5700 5.5500 1.6700 ;
      RECT 3.4200 1.3900 3.5900 1.4800 ;
      RECT 3.5000 0.5700 3.5900 1.3900 ;
      RECT 1.7300 0.5700 1.8200 1.2200 ;
      RECT 1.6750 1.2200 1.8200 1.4100 ;
      RECT 1.8750 1.8300 6.1200 1.9200 ;
      RECT 6.0300 1.4950 6.1200 1.8300 ;
      RECT 6.0300 1.4050 6.1300 1.4950 ;
      RECT 6.0400 0.8850 6.1300 1.4050 ;
      RECT 6.0300 0.7950 6.1300 0.8850 ;
      RECT 6.0300 0.6750 6.1200 0.7950 ;
      RECT 3.1550 1.9200 3.3250 1.9900 ;
  END
END SDFFSQN_X2M_A12TH

MACRO SDFFSQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7400 ;
        RECT 1.0300 0.3200 1.1300 0.6200 ;
        RECT 3.9700 0.3200 4.3400 0.3800 ;
        RECT 6.1500 0.3200 6.2500 0.4950 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3800 1.2100 1.5500 1.4000 ;
        RECT 1.3800 1.0400 1.4800 1.2100 ;
    END
    ANTENNAGATEAREA 0.0954 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 6.0950 2.0300 6.2650 2.0800 ;
        RECT 3.9050 2.0200 4.0750 2.0800 ;
        RECT 1.0050 1.8000 1.1050 2.0800 ;
        RECT 0.0750 1.7250 0.1750 2.0800 ;
    END
  END VDD

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1000 1.0100 1.3900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2500 0.7250 6.3500 1.1450 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0950 1.2500 5.7150 1.3500 ;
        RECT 5.0950 1.3500 5.1950 1.7200 ;
        RECT 5.6150 1.3500 5.7150 1.7300 ;
        RECT 5.6150 0.8300 5.7150 1.2500 ;
        RECT 5.0600 0.7300 5.7150 0.8300 ;
    END
    ANTENNADIFFAREA 0.5598 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8200 1.0300 2.9700 1.4150 ;
    END
    ANTENNAGATEAREA 0.1134 ;
  END SN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.3350 1.8200 0.7500 1.9200 ;
      RECT 0.3350 0.5300 0.4350 1.8200 ;
      RECT 0.3350 0.4300 0.7350 0.5300 ;
      RECT 1.4650 1.6100 1.5650 1.9600 ;
      RECT 0.5250 1.5200 1.5650 1.6100 ;
      RECT 0.5250 0.7950 1.5900 0.8850 ;
      RECT 1.4900 0.4900 1.5900 0.7950 ;
      RECT 0.5250 0.8850 0.6250 1.5200 ;
      RECT 1.6950 1.6350 1.9650 1.7250 ;
      RECT 1.8750 0.9400 1.9650 1.6350 ;
      RECT 1.8750 0.8500 2.6800 0.9400 ;
      RECT 2.5900 0.9400 2.6800 1.3250 ;
      RECT 2.2550 1.6150 3.1950 1.7150 ;
      RECT 3.0950 0.7600 3.1950 1.6150 ;
      RECT 2.9350 0.6600 3.1950 0.7600 ;
      RECT 2.2550 1.1800 2.3550 1.6150 ;
      RECT 3.3100 1.4650 4.3950 1.5550 ;
      RECT 4.3050 1.1800 4.3950 1.4650 ;
      RECT 3.3100 0.7850 3.4000 1.4650 ;
      RECT 4.3050 1.0900 4.7800 1.1800 ;
      RECT 4.4950 1.3700 4.9700 1.4700 ;
      RECT 4.8700 0.9050 4.9700 1.3700 ;
      RECT 3.8050 0.8050 4.9700 0.9050 ;
      RECT 3.8050 0.9050 3.9050 1.3650 ;
      RECT 2.7300 0.4800 5.9600 0.5700 ;
      RECT 5.8700 0.5700 5.9600 1.7400 ;
      RECT 1.6800 0.6000 2.8200 0.6900 ;
      RECT 2.7300 0.5700 2.8200 0.6000 ;
      RECT 3.5150 0.5700 3.6150 1.3700 ;
      RECT 1.6400 1.2450 1.7700 1.4150 ;
      RECT 1.6800 0.6900 1.7700 1.2450 ;
      RECT 1.8200 1.8300 6.5550 1.9200 ;
      RECT 6.4550 1.5000 6.5550 1.8300 ;
      RECT 6.0550 1.4100 6.5550 1.5000 ;
      RECT 6.4550 0.5650 6.5550 1.4100 ;
      RECT 6.3750 0.4650 6.5550 0.5650 ;
      RECT 6.0550 1.2900 6.1450 1.4100 ;
      RECT 3.4700 1.9200 3.6400 1.9750 ;
      RECT 1.8200 1.9200 1.9900 1.9600 ;
  END
END SDFFSQN_X3M_A12TH

MACRO SDFFSQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.9150 ;
        RECT 1.0900 0.3200 1.2600 0.6900 ;
        RECT 2.5700 0.3200 2.7400 0.7200 ;
        RECT 5.6900 0.3200 5.7900 0.9000 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0600 0.1700 1.5450 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0200 1.0100 1.1500 1.3500 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 4.7400 1.9700 4.9500 2.0800 ;
        RECT 5.6150 1.9700 5.8250 2.0800 ;
        RECT 0.0800 1.7000 0.1800 2.0800 ;
        RECT 1.0900 1.6600 1.2600 2.0800 ;
    END
  END VDD

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.1900 3.0550 1.3600 ;
        RECT 2.8500 1.3600 2.9500 1.4600 ;
        RECT 2.8500 1.0150 2.9500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END SN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.7200 5.1900 1.6500 ;
    END
    ANTENNADIFFAREA 0.1358 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.0350 1.5650 1.3900 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.0100 5.8000 1.4050 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3450 1.7400 0.8300 1.8300 ;
      RECT 0.3450 0.6000 0.4350 1.7400 ;
      RECT 0.3450 0.5100 0.6500 0.6000 ;
      RECT 0.5450 1.4800 1.7100 1.5700 ;
      RECT 0.5450 0.7800 1.7100 0.8700 ;
      RECT 0.5450 0.8700 0.6450 1.4800 ;
      RECT 1.8000 1.5100 2.0800 1.6000 ;
      RECT 1.9900 1.0800 2.0800 1.5100 ;
      RECT 1.9900 0.9900 2.7300 1.0800 ;
      RECT 2.6400 1.0800 2.7300 1.3050 ;
      RECT 1.9900 0.8600 2.0800 0.9900 ;
      RECT 1.9900 0.7600 2.1800 0.8600 ;
      RECT 2.3000 1.5800 3.2700 1.6700 ;
      RECT 3.1800 0.9800 3.2700 1.5800 ;
      RECT 3.0850 0.8900 3.2700 0.9800 ;
      RECT 3.0850 0.7050 3.1750 0.8900 ;
      RECT 2.3000 1.1850 2.3900 1.5800 ;
      RECT 3.3900 1.5400 4.4000 1.6300 ;
      RECT 4.3100 1.1750 4.4000 1.5400 ;
      RECT 3.3900 0.7050 3.4800 1.5400 ;
      RECT 4.3100 1.0850 4.7500 1.1750 ;
      RECT 4.5150 1.3750 4.6050 1.6550 ;
      RECT 4.5150 1.2850 4.9400 1.3750 ;
      RECT 4.8500 0.8550 4.9400 1.2850 ;
      RECT 3.8300 0.7650 4.9400 0.8550 ;
      RECT 3.8300 0.8550 3.9200 1.3950 ;
      RECT 2.8500 0.4900 5.4500 0.5800 ;
      RECT 5.3600 0.5800 5.4500 1.4500 ;
      RECT 2.3700 0.8100 2.9400 0.9000 ;
      RECT 2.8500 0.5800 2.9400 0.8100 ;
      RECT 3.6000 0.5800 3.6900 1.4050 ;
      RECT 3.2300 0.4800 3.4000 0.4900 ;
      RECT 1.6950 1.2350 1.8900 1.3250 ;
      RECT 1.8000 0.6200 1.8900 1.2350 ;
      RECT 1.8000 0.5300 2.4600 0.6200 ;
      RECT 2.3700 0.6200 2.4600 0.8100 ;
      RECT 1.8850 1.7900 6.1050 1.8800 ;
      RECT 6.0150 0.7050 6.1050 1.7900 ;
  END
END SDFFSQ_X0P5M_A12TH

MACRO SDFFSQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.9200 ;
        RECT 1.0950 0.3200 1.2650 0.7400 ;
        RECT 2.5600 0.3200 2.7300 0.5400 ;
        RECT 4.1650 0.3200 4.3750 0.5350 ;
        RECT 4.8250 0.3200 4.9950 0.3700 ;
        RECT 5.6950 0.3200 5.7850 0.9200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.8100 2.0400 3.0200 2.0800 ;
        RECT 1.1250 1.9150 1.2350 2.0800 ;
        RECT 0.0850 1.6800 0.1850 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.2200 1.6700 ;
        RECT 5.1200 0.7850 5.2200 1.4100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.1650 5.7500 1.4950 ;
        RECT 5.6500 1.0750 5.9050 1.1650 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1700 1.5050 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0300 1.0600 1.1500 1.4500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4300 1.0800 1.5700 1.4900 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8450 1.1850 3.0450 1.4100 ;
    END
    ANTENNAGATEAREA 0.0792 ;
  END SN
  OBS
    LAYER M1 ;
      RECT 0.3450 1.8800 0.7650 1.9700 ;
      RECT 0.3450 0.5900 0.4450 1.8800 ;
      RECT 0.3450 0.4900 0.6700 0.5900 ;
      RECT 0.5950 1.6800 1.7150 1.7700 ;
      RECT 0.5550 0.8300 1.6750 0.9200 ;
      RECT 1.5850 0.5100 1.6750 0.8300 ;
      RECT 0.5950 0.9200 0.6850 1.6800 ;
      RECT 1.8050 1.6250 2.0800 1.7150 ;
      RECT 1.9900 1.1700 2.0800 1.6250 ;
      RECT 1.9900 1.0800 2.7500 1.1700 ;
      RECT 2.6600 1.1700 2.7500 1.2900 ;
      RECT 1.9900 0.7450 2.0800 1.0800 ;
      RECT 2.2500 1.6300 3.2350 1.7300 ;
      RECT 3.1350 0.7550 3.2350 1.6300 ;
      RECT 2.2500 1.2900 2.3500 1.6300 ;
      RECT 3.3750 1.6500 4.3750 1.7400 ;
      RECT 4.2850 1.1700 4.3750 1.6500 ;
      RECT 3.3750 0.9650 3.4650 1.6500 ;
      RECT 4.2850 1.0800 4.7400 1.1700 ;
      RECT 3.3750 0.7550 3.5000 0.9650 ;
      RECT 4.5350 1.4150 4.6250 1.7400 ;
      RECT 4.5350 1.3250 4.9600 1.4150 ;
      RECT 4.8700 0.9350 4.9600 1.3250 ;
      RECT 3.8200 0.8450 4.9600 0.9350 ;
      RECT 3.8200 0.9350 3.9100 1.5350 ;
      RECT 3.5900 0.6350 5.4800 0.6600 ;
      RECT 5.3900 0.6600 5.4800 1.6550 ;
      RECT 4.6150 0.5700 5.4800 0.6350 ;
      RECT 3.5900 0.6600 4.7050 0.7250 ;
      RECT 1.6800 1.3500 1.8700 1.4400 ;
      RECT 1.7800 0.6050 1.8700 1.3500 ;
      RECT 1.7800 0.5150 2.4400 0.6050 ;
      RECT 2.3500 0.6050 2.4400 0.6300 ;
      RECT 2.3500 0.6300 2.9400 0.7200 ;
      RECT 2.8500 0.5700 2.9400 0.6300 ;
      RECT 2.8500 0.4800 3.6800 0.5700 ;
      RECT 3.5900 0.5700 3.6800 0.6350 ;
      RECT 3.2650 0.4350 3.4750 0.4800 ;
      RECT 3.5900 0.7250 3.6800 1.5400 ;
      RECT 1.9150 1.8300 6.1200 1.9200 ;
      RECT 6.0300 0.7450 6.1200 1.8300 ;
      RECT 3.2350 1.9200 3.4450 1.9850 ;
      RECT 1.9150 1.9200 2.1250 1.9600 ;
  END
END SDFFSQ_X1M_A12TH

MACRO SDFFSQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9000 ;
        RECT 1.0750 0.3200 1.1950 0.6400 ;
        RECT 2.5250 0.3200 2.6250 0.4650 ;
        RECT 5.7150 0.3200 5.8150 0.8900 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9850 1.4100 5.1500 1.6700 ;
        RECT 4.9850 0.7100 5.0850 1.4100 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0900 2.9700 1.5100 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END SN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8200 1.0100 5.9500 1.3350 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 4.6900 2.0400 4.8600 2.0800 ;
        RECT 5.2100 2.0400 5.3800 2.0800 ;
        RECT 5.7000 2.0400 5.8700 2.0800 ;
        RECT 2.7300 2.0100 2.9400 2.0800 ;
        RECT 1.0700 1.8250 1.1600 2.0800 ;
        RECT 0.0800 1.7000 0.1700 2.0800 ;
    END
  END VDD

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2900 0.9500 1.4900 ;
        RECT 0.8500 1.1200 1.0350 1.2900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 1.0650 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0792 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8300 0.8050 1.9200 ;
      RECT 0.3400 0.5500 0.4300 1.8300 ;
      RECT 0.3400 0.4600 0.6150 0.5500 ;
      RECT 1.5300 1.7050 1.6200 1.9850 ;
      RECT 0.5700 1.6150 1.6200 1.7050 ;
      RECT 0.5700 0.7800 1.6300 0.8700 ;
      RECT 1.5400 0.4750 1.6300 0.7800 ;
      RECT 0.5700 0.8700 0.6600 1.6150 ;
      RECT 1.7300 1.5700 2.0300 1.6600 ;
      RECT 1.9400 0.9100 2.0300 1.5700 ;
      RECT 1.9400 0.8200 2.7250 0.9100 ;
      RECT 2.6350 0.9100 2.7250 1.2900 ;
      RECT 2.2200 1.6500 3.1500 1.7400 ;
      RECT 3.0600 0.8800 3.1500 1.6500 ;
      RECT 2.9250 0.7900 3.1500 0.8800 ;
      RECT 2.2200 1.2650 2.3100 1.6500 ;
      RECT 3.2600 1.6500 4.2550 1.7400 ;
      RECT 3.2600 1.5950 3.4550 1.6500 ;
      RECT 4.1650 1.1700 4.2550 1.6500 ;
      RECT 3.2600 0.7600 3.3500 1.5950 ;
      RECT 4.1650 1.0800 4.5700 1.1700 ;
      RECT 4.4150 1.4150 4.5050 1.6950 ;
      RECT 4.4150 1.3250 4.8850 1.4150 ;
      RECT 4.7950 0.8750 4.8850 1.3250 ;
      RECT 3.7100 0.7850 4.8850 0.8750 ;
      RECT 3.7100 0.8750 3.8000 1.4950 ;
      RECT 2.9500 0.4800 5.5450 0.5700 ;
      RECT 5.4550 0.5700 5.5450 1.6700 ;
      RECT 3.4400 1.3900 3.6100 1.4800 ;
      RECT 3.5200 0.5700 3.6100 1.3900 ;
      RECT 2.9500 0.5700 3.0400 0.5750 ;
      RECT 3.3350 0.4100 3.5450 0.4800 ;
      RECT 1.7250 0.5750 3.0400 0.6650 ;
      RECT 1.7250 0.6650 1.8150 1.2200 ;
      RECT 1.6750 1.2200 1.8150 1.4100 ;
      RECT 1.8750 1.8300 5.9450 1.9200 ;
      RECT 5.8550 1.5350 5.9450 1.8300 ;
      RECT 5.8550 1.4450 6.1550 1.5350 ;
      RECT 6.0650 0.8350 6.1550 1.4450 ;
      RECT 5.9650 0.7450 6.1550 0.8350 ;
      RECT 3.1550 1.9200 3.3650 1.9900 ;
  END
END SDFFSQ_X2M_A12TH

MACRO SDFFSQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.9200 ;
        RECT 1.0850 0.3200 1.1850 0.6100 ;
        RECT 2.5600 0.3200 2.6600 0.5600 ;
        RECT 4.7650 0.3200 4.9350 0.5200 ;
        RECT 5.3250 0.3200 5.4150 0.4600 ;
        RECT 6.1450 0.3200 6.2450 0.7150 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 3.9300 2.0200 4.1400 2.0800 ;
        RECT 2.7650 2.0100 2.9750 2.0800 ;
        RECT 6.1400 1.8600 6.2400 2.0800 ;
        RECT 1.0850 1.8000 1.1850 2.0800 ;
        RECT 0.0850 1.6800 0.1850 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.0400 1.5650 1.3900 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.0100 1.1500 1.3150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.9650 6.2950 1.1350 ;
        RECT 6.0500 1.1350 6.1500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0600 1.2500 5.7150 1.3500 ;
        RECT 5.0600 1.3500 5.1600 1.6900 ;
        RECT 5.5850 1.3500 5.7150 1.6700 ;
        RECT 5.5800 0.9100 5.7150 1.2500 ;
        RECT 5.0250 0.8100 5.7150 0.9100 ;
    END
    ANTENNADIFFAREA 0.571425 ;
  END Q

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0300 3.0100 1.4150 ;
    END
    ANTENNAGATEAREA 0.1068 ;
  END SN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.075 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.3450 1.7750 0.7850 1.8750 ;
      RECT 0.3450 0.5950 0.4450 1.7750 ;
      RECT 0.3450 0.4950 0.6350 0.5950 ;
      RECT 1.5450 1.6000 1.6450 1.9200 ;
      RECT 0.5400 1.5100 1.6450 1.6000 ;
      RECT 0.5400 0.8300 1.6500 0.9200 ;
      RECT 1.5600 0.4900 1.6500 0.8300 ;
      RECT 0.5400 0.9200 0.6300 1.5100 ;
      RECT 1.7600 1.4950 2.0400 1.5850 ;
      RECT 1.9500 0.9200 2.0400 1.4950 ;
      RECT 1.9500 0.8300 2.7200 0.9200 ;
      RECT 2.6300 0.9200 2.7200 1.2400 ;
      RECT 2.2800 1.6100 3.2350 1.7100 ;
      RECT 3.1350 0.8050 3.2350 1.6100 ;
      RECT 2.9700 0.7050 3.2350 0.8050 ;
      RECT 2.2800 1.1800 2.3800 1.6100 ;
      RECT 3.3500 1.4650 4.4350 1.5550 ;
      RECT 4.3450 1.1600 4.4350 1.4650 ;
      RECT 3.3500 0.7850 3.4400 1.4650 ;
      RECT 4.3450 1.0600 4.7400 1.1600 ;
      RECT 4.8350 1.0500 5.3400 1.1500 ;
      RECT 4.5400 1.3750 4.6400 1.6700 ;
      RECT 4.5400 1.2750 4.9250 1.3750 ;
      RECT 4.8350 1.1500 4.9250 1.2750 ;
      RECT 4.8350 0.9250 4.9250 1.0500 ;
      RECT 3.8600 0.8250 4.9250 0.9250 ;
      RECT 3.8600 0.9250 3.9600 1.3650 ;
      RECT 3.5750 0.6100 5.9550 0.7000 ;
      RECT 5.8650 0.7000 5.9550 1.5000 ;
      RECT 1.7400 0.7400 1.8300 1.4050 ;
      RECT 2.0300 0.5950 2.2400 0.6500 ;
      RECT 1.7400 0.6500 2.8600 0.7400 ;
      RECT 2.7700 0.5700 2.8600 0.6500 ;
      RECT 2.7700 0.4800 3.6650 0.5700 ;
      RECT 3.5750 0.5700 3.6650 0.6100 ;
      RECT 3.5750 0.7000 3.6650 1.3700 ;
      RECT 5.8850 1.6550 6.5050 1.7450 ;
      RECT 6.4150 0.4600 6.5050 1.6550 ;
      RECT 3.4900 1.9200 3.7000 1.9750 ;
      RECT 1.8850 1.8300 5.9750 1.9200 ;
      RECT 5.8850 1.7450 5.9750 1.8300 ;
  END
END SDFFSQ_X3M_A12TH

MACRO SDFFSQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.9200 ;
        RECT 1.1250 0.3200 1.2150 0.6100 ;
        RECT 6.7500 0.3200 6.8500 0.9050 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 2.8100 2.0250 2.9800 2.0800 ;
        RECT 1.1050 1.8200 1.2050 2.0800 ;
        RECT 6.7050 1.7900 6.7950 2.0800 ;
        RECT 0.0850 1.6800 0.1850 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 1.3500 5.9700 1.6500 ;
        RECT 5.3500 1.2500 5.9700 1.3500 ;
        RECT 5.3500 1.3500 5.4500 1.6700 ;
        RECT 5.8700 0.8200 5.9700 1.2500 ;
        RECT 5.2900 0.7200 5.9700 0.8200 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 1.1650 6.7500 1.4000 ;
        RECT 6.6500 1.0750 6.9250 1.1650 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1700 1.5050 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8300 1.2100 3.0350 1.3900 ;
        RECT 2.8300 0.7500 2.9200 1.2100 ;
        RECT 2.8300 0.6600 3.4000 0.7500 ;
        RECT 3.3100 0.7500 3.4000 1.6500 ;
        RECT 3.3100 1.6500 4.4500 1.7400 ;
    END
    ANTENNAGATEAREA 0.1044 ;
  END SN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.0200 1.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4300 1.0600 1.5700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3500 1.7800 0.8150 1.8700 ;
      RECT 0.3500 0.5400 0.4400 1.7800 ;
      RECT 0.3500 0.4500 0.6550 0.5400 ;
      RECT 1.5650 1.6050 1.6650 1.9300 ;
      RECT 0.5700 1.5150 1.6650 1.6050 ;
      RECT 0.5700 0.8100 1.6750 0.9000 ;
      RECT 1.5850 0.5100 1.6750 0.8100 ;
      RECT 0.5700 0.9250 0.6600 1.5150 ;
      RECT 0.5700 0.9000 0.7500 0.9250 ;
      RECT 1.7900 1.5450 2.0850 1.6350 ;
      RECT 1.9950 0.9400 2.0850 1.5450 ;
      RECT 1.9950 0.8500 2.7200 0.9400 ;
      RECT 2.6300 0.9400 2.7200 1.3500 ;
      RECT 2.2850 1.6400 3.2200 1.7300 ;
      RECT 3.1300 0.9550 3.2200 1.6400 ;
      RECT 3.0100 0.8650 3.2200 0.9550 ;
      RECT 2.2850 1.2100 2.3750 1.6400 ;
      RECT 3.4950 1.4600 4.4950 1.5500 ;
      RECT 4.4050 1.1700 4.4950 1.4600 ;
      RECT 3.4950 0.7350 3.5850 1.4600 ;
      RECT 4.4050 1.0800 4.9550 1.1700 ;
      RECT 5.0800 1.0500 5.7100 1.1400 ;
      RECT 4.7750 1.6300 5.1700 1.7200 ;
      RECT 5.0800 1.1400 5.1700 1.6300 ;
      RECT 5.0800 0.8500 5.1700 1.0500 ;
      RECT 3.9450 0.7600 5.1700 0.8500 ;
      RECT 3.9450 0.8500 4.0350 1.3600 ;
      RECT 2.2600 0.4800 6.5350 0.5700 ;
      RECT 6.4450 0.5700 6.5350 1.4700 ;
      RECT 3.7000 0.5700 3.7900 1.3700 ;
      RECT 1.6850 1.2700 1.8900 1.3600 ;
      RECT 1.8000 0.6800 1.8900 1.2700 ;
      RECT 1.8000 0.5900 2.3500 0.6800 ;
      RECT 2.2600 0.5700 2.3500 0.5900 ;
      RECT 6.2450 1.6100 7.1050 1.7000 ;
      RECT 7.0150 0.5800 7.1050 1.6100 ;
      RECT 1.9250 1.8300 6.3450 1.9200 ;
      RECT 6.2450 1.7000 6.3450 1.8300 ;
      RECT 6.2450 1.0050 6.3450 1.6100 ;
      RECT 3.6350 1.9200 3.8050 1.9900 ;
  END
END SDFFSQ_X4M_A12TH

MACRO SDFFSRPQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.0650 0.3200 0.1850 0.4100 ;
        RECT 1.0150 0.3200 1.1150 0.7200 ;
        RECT 3.8250 0.3200 4.1150 0.3850 ;
        RECT 5.8300 0.3200 6.0000 0.3850 ;
        RECT 6.6750 0.3200 6.8450 0.7400 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4100 1.4600 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0950 4.2400 1.2650 ;
        RECT 4.0500 0.8550 4.1800 1.0950 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1850 1.2050 5.3550 1.4650 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.8500 6.1500 1.5850 ;
        RECT 6.0500 1.5850 6.2950 1.6850 ;
        RECT 6.0500 0.7500 6.3000 0.8500 ;
    END
    ANTENNADIFFAREA 0.217775 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 2.0900 2.0600 2.4600 2.0800 ;
        RECT 3.1150 2.0400 3.5200 2.0800 ;
        RECT 3.6800 2.0400 4.0500 2.0800 ;
        RECT 6.7050 2.0300 7.0750 2.0800 ;
        RECT 5.8300 2.0200 6.0000 2.0800 ;
        RECT 1.0050 1.9000 1.1250 2.0800 ;
        RECT 3.1150 2.0350 3.3250 2.0400 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4200 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0150 0.9600 1.4850 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 1.1550 6.7500 1.3900 ;
        RECT 6.6500 1.0450 6.9200 1.1550 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3150 1.8800 0.7300 1.9700 ;
      RECT 0.3150 1.7900 0.4050 1.8800 ;
      RECT 0.0600 1.7000 0.4050 1.7900 ;
      RECT 0.0600 0.5000 0.6900 0.5900 ;
      RECT 0.6000 0.4100 0.7900 0.5000 ;
      RECT 0.0600 0.5900 0.1500 1.7000 ;
      RECT 1.0700 1.6000 1.6750 1.7000 ;
      RECT 0.4450 0.8100 1.6350 0.9000 ;
      RECT 1.5450 0.7150 1.6350 0.8100 ;
      RECT 0.4950 1.7000 1.1600 1.7900 ;
      RECT 1.0700 0.9000 1.1600 1.6000 ;
      RECT 0.4950 1.5450 0.5850 1.7000 ;
      RECT 0.4450 0.9000 0.6150 0.9100 ;
      RECT 1.7800 1.6000 1.9950 1.6900 ;
      RECT 1.9050 1.1900 1.9950 1.6000 ;
      RECT 1.9050 1.1000 2.9100 1.1900 ;
      RECT 2.8200 1.1900 2.9100 1.2900 ;
      RECT 1.9050 0.6800 1.9950 1.1000 ;
      RECT 2.7350 0.7800 2.8250 0.9150 ;
      RECT 2.7350 0.6900 3.3450 0.7800 ;
      RECT 3.2550 0.7800 3.3450 0.9150 ;
      RECT 2.6650 1.4700 2.7550 1.7400 ;
      RECT 2.2100 1.3800 3.6300 1.4700 ;
      RECT 2.2100 1.3000 2.3000 1.3800 ;
      RECT 3.5400 1.1000 3.6300 1.3800 ;
      RECT 3.0350 1.0100 3.6300 1.1000 ;
      RECT 3.0350 0.9600 3.1250 1.0100 ;
      RECT 3.5300 0.7250 3.6300 1.0100 ;
      RECT 2.9550 0.8700 3.1250 0.9600 ;
      RECT 4.5600 0.6600 5.5300 0.7500 ;
      RECT 5.4400 0.7500 5.5300 0.9450 ;
      RECT 5.4400 0.9450 5.6000 1.1150 ;
      RECT 3.7950 1.6450 4.6500 1.7350 ;
      RECT 4.5600 0.7500 4.6500 1.6450 ;
      RECT 3.7950 1.5100 3.8850 1.6450 ;
      RECT 3.7600 1.3400 3.8850 1.5100 ;
      RECT 3.7950 0.7250 3.8850 1.3400 ;
      RECT 4.9400 1.6400 5.9000 1.7300 ;
      RECT 5.8100 0.7700 5.9000 1.6400 ;
      RECT 5.6250 0.6800 5.9000 0.7700 ;
      RECT 4.9400 1.3500 5.0300 1.6400 ;
      RECT 1.7250 0.4800 6.5150 0.5700 ;
      RECT 6.4250 0.5700 6.5150 1.7400 ;
      RECT 4.3600 0.5700 4.4500 1.5350 ;
      RECT 1.7250 0.5700 1.8150 1.4550 ;
      RECT 1.8950 1.8300 7.1050 1.9200 ;
      RECT 7.0150 0.5600 7.1050 1.8300 ;
      RECT 4.7500 0.8850 4.8400 1.8300 ;
  END
END SDFFSRPQ_X0P5M_A12TH

MACRO SDFFSRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.0750 0.3200 0.2150 0.4650 ;
        RECT 1.0350 0.3200 1.1350 0.7200 ;
        RECT 3.7750 0.3200 4.1850 0.3700 ;
        RECT 5.3750 0.3200 5.4950 0.3500 ;
        RECT 5.6350 0.3200 6.0450 0.3350 ;
        RECT 6.6800 0.3200 6.8500 0.8500 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4100 1.5050 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0950 4.2500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1800 1.0100 5.3500 1.3150 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 1.2900 6.2450 1.6600 ;
        RECT 6.0500 0.8850 6.1500 1.2900 ;
        RECT 6.0500 0.7150 6.2850 0.8850 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 5.6550 2.0600 6.0450 2.0800 ;
        RECT 2.1550 2.0300 2.5650 2.0800 ;
        RECT 3.1150 2.0300 3.5250 2.0800 ;
        RECT 3.7150 2.0300 4.1200 2.0800 ;
        RECT 1.0000 1.8800 1.1700 2.0800 ;
        RECT 6.6850 1.8200 6.8550 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9600 1.5100 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 1.0100 6.9050 1.1900 ;
        RECT 6.6500 1.1900 6.7700 1.5050 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3350 1.8800 0.7500 1.9700 ;
      RECT 0.3350 1.7900 0.4250 1.8800 ;
      RECT 0.0600 1.7000 0.4250 1.7900 ;
      RECT 0.0600 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5200 0.5100 0.6000 ;
      RECT 0.4200 0.4300 0.8100 0.5200 ;
      RECT 0.0600 0.6900 0.1500 1.7000 ;
      RECT 0.5150 1.7000 1.6300 1.7900 ;
      RECT 0.4650 0.8100 1.5900 0.9000 ;
      RECT 1.5000 0.6900 1.5900 0.8100 ;
      RECT 1.0700 0.9000 1.1600 1.7000 ;
      RECT 0.5150 1.5350 0.6050 1.7000 ;
      RECT 0.4650 0.9000 0.6350 0.9300 ;
      RECT 1.7250 1.5900 1.9500 1.6800 ;
      RECT 1.8600 1.1900 1.9500 1.5900 ;
      RECT 1.8600 1.1000 2.9200 1.1900 ;
      RECT 2.8300 1.1900 2.9200 1.4600 ;
      RECT 1.8600 0.6800 1.9500 1.1000 ;
      RECT 2.6700 0.6700 3.3800 0.7600 ;
      RECT 2.1550 1.6200 3.6050 1.7100 ;
      RECT 3.4800 1.5050 3.6050 1.6200 ;
      RECT 2.1550 1.3050 2.2450 1.6200 ;
      RECT 3.5150 0.9600 3.6050 1.5050 ;
      RECT 2.9300 0.8700 3.6050 0.9600 ;
      RECT 3.5150 0.7550 3.6050 0.8700 ;
      RECT 4.5900 0.6700 5.5900 0.7600 ;
      RECT 5.5000 0.7600 5.5900 1.0400 ;
      RECT 5.5000 1.0400 5.6100 1.2100 ;
      RECT 3.7400 1.6450 4.6800 1.7350 ;
      RECT 4.5900 0.7600 4.6800 1.6450 ;
      RECT 3.7400 1.4950 3.8800 1.6450 ;
      RECT 3.7900 0.7550 3.8800 1.4950 ;
      RECT 4.9800 1.6400 5.8500 1.7300 ;
      RECT 5.7600 1.1950 5.8500 1.6400 ;
      RECT 5.7600 1.0250 5.8900 1.1950 ;
      RECT 5.7600 0.8850 5.8500 1.0250 ;
      RECT 5.6800 0.6950 5.8500 0.8850 ;
      RECT 4.9800 1.3700 5.0700 1.6400 ;
      RECT 6.3950 1.3600 6.5300 1.5500 ;
      RECT 6.3950 0.8700 6.4850 1.3600 ;
      RECT 6.3950 0.7000 6.5250 0.8700 ;
      RECT 6.3950 0.5700 6.4850 0.7000 ;
      RECT 1.6800 0.4800 6.4850 0.5700 ;
      RECT 4.4000 0.5700 4.4900 1.5350 ;
      RECT 1.6800 0.5700 1.7700 1.2850 ;
      RECT 1.9250 0.4600 2.0950 0.4800 ;
      RECT 1.6600 1.2850 1.7700 1.4550 ;
      RECT 6.4500 1.6400 7.1050 1.7300 ;
      RECT 7.0150 0.6600 7.1050 1.6400 ;
      RECT 1.8650 1.8300 6.5400 1.9200 ;
      RECT 6.4500 1.7300 6.5400 1.8300 ;
      RECT 4.7900 0.8850 4.8800 1.8300 ;
  END
END SDFFSRPQ_X1M_A12TH

MACRO SDFFSRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.4450 0.3200 ;
        RECT 0.0750 0.3200 0.2150 0.4650 ;
        RECT 1.0350 0.3200 1.1350 0.7200 ;
        RECT 3.9750 0.3200 4.1450 0.3500 ;
        RECT 6.8250 0.3200 6.9950 0.7600 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4100 1.4600 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0450 1.1600 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.1224 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1650 1.0100 5.3500 1.1900 ;
        RECT 5.1650 1.1900 5.2550 1.3400 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 1.2900 6.2050 1.6600 ;
        RECT 6.0500 0.8850 6.1500 1.2900 ;
        RECT 6.0500 0.7150 6.2450 0.8850 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.4450 2.7200 ;
        RECT 3.1150 2.0650 3.5250 2.0800 ;
        RECT 2.1550 2.0550 2.5650 2.0800 ;
        RECT 5.8400 2.0400 5.9800 2.0800 ;
        RECT 5.3650 2.0350 5.5050 2.0800 ;
        RECT 3.8900 2.0300 4.0950 2.0800 ;
        RECT 1.0250 1.9350 1.1450 2.0800 ;
        RECT 6.8300 1.8100 7.0000 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9700 1.4650 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8500 1.1600 6.9500 1.3900 ;
        RECT 6.8500 1.0500 7.0700 1.1600 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 6.6050 1.6300 7.2750 1.7200 ;
      RECT 7.1600 1.4450 7.2750 1.6300 ;
      RECT 7.1850 0.7950 7.2750 1.4450 ;
      RECT 7.1600 0.6250 7.2750 0.7950 ;
      RECT 6.5250 1.9200 6.6950 1.9500 ;
      RECT 1.8650 1.8300 6.6950 1.9200 ;
      RECT 6.6050 1.7200 6.6950 1.8300 ;
      RECT 4.7650 0.8850 4.8550 1.8300 ;
      RECT 3.2450 1.2450 3.3350 1.8300 ;
      RECT 3.2450 1.0750 3.4250 1.2450 ;
      RECT 0.3350 1.8800 0.7500 1.9700 ;
      RECT 0.3350 1.7900 0.4250 1.8800 ;
      RECT 0.0600 1.7000 0.4250 1.7900 ;
      RECT 0.0600 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5200 0.5100 0.6000 ;
      RECT 0.4200 0.4300 0.8100 0.5200 ;
      RECT 0.0600 0.6900 0.1500 1.7000 ;
      RECT 0.5150 1.7000 1.6300 1.7900 ;
      RECT 0.4650 0.8100 1.5900 0.9000 ;
      RECT 1.5000 0.4900 1.5900 0.8100 ;
      RECT 1.0700 0.9000 1.1600 1.7000 ;
      RECT 0.5150 1.5350 0.6050 1.7000 ;
      RECT 0.4650 0.9000 0.6350 0.9300 ;
      RECT 1.7250 1.5900 1.9500 1.6800 ;
      RECT 1.8600 1.1750 1.9500 1.5900 ;
      RECT 1.8600 1.0850 2.9200 1.1750 ;
      RECT 2.8300 1.1750 2.9200 1.2800 ;
      RECT 1.8600 0.6800 1.9500 1.0850 ;
      RECT 2.6700 0.6700 3.4000 0.7600 ;
      RECT 3.4350 1.5400 3.6050 1.7100 ;
      RECT 3.5150 0.9600 3.6050 1.5400 ;
      RECT 2.9300 0.8700 3.6050 0.9600 ;
      RECT 3.0450 0.9600 3.1350 1.4400 ;
      RECT 3.5150 0.7350 3.6050 0.8700 ;
      RECT 2.1850 1.4400 3.1350 1.5300 ;
      RECT 2.1850 1.2850 2.2750 1.4400 ;
      RECT 4.5650 0.6600 5.5600 0.7500 ;
      RECT 5.4700 0.7500 5.5600 1.1100 ;
      RECT 5.4700 1.1100 5.5850 1.2800 ;
      RECT 3.6950 1.6450 4.6550 1.7350 ;
      RECT 4.5650 0.7500 4.6550 1.6450 ;
      RECT 3.6950 0.9100 3.7850 1.6450 ;
      RECT 3.6950 0.7300 3.8800 0.9100 ;
      RECT 4.9550 1.6400 5.8450 1.7300 ;
      RECT 5.7550 0.9500 5.8450 1.6400 ;
      RECT 5.6500 0.7350 5.8450 0.9500 ;
      RECT 4.9550 1.3500 5.0450 1.6400 ;
      RECT 1.6800 0.4800 6.6700 0.5700 ;
      RECT 6.5800 0.5700 6.6700 1.5400 ;
      RECT 4.0150 0.5700 4.1050 1.0000 ;
      RECT 4.3750 0.5700 4.4650 1.5350 ;
      RECT 1.6600 1.2850 1.7700 1.4550 ;
      RECT 1.6800 0.5700 1.7700 1.2850 ;
      RECT 1.9250 0.4550 2.0950 0.4800 ;
  END
END SDFFSRPQ_X2M_A12TH

MACRO SDFFSRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.0750 0.3200 0.2150 0.4650 ;
        RECT 1.0350 0.3200 1.1350 0.6700 ;
        RECT 3.9250 0.3200 4.1350 0.3700 ;
        RECT 5.2600 0.3200 5.4700 0.3600 ;
        RECT 5.7700 0.3200 5.8900 0.3900 ;
        RECT 6.2500 0.3200 6.4500 0.3700 ;
        RECT 7.0600 0.3200 7.2300 0.6900 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4100 1.4600 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0050 1.0450 5.2650 1.1550 ;
        RECT 5.1550 0.8700 5.2650 1.0450 ;
    END
    ANTENNAGATEAREA 0.1254 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0200 1.0500 3.1500 1.4100 ;
    END
    ANTENNAGATEAREA 0.1134 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0050 0.8500 6.6550 0.9500 ;
        RECT 6.4500 0.9500 6.5500 1.2900 ;
        RECT 6.0050 0.7050 6.1750 0.8500 ;
        RECT 6.5650 0.7050 6.6550 0.8500 ;
        RECT 6.0400 1.2900 6.6550 1.3900 ;
        RECT 6.0400 1.3900 6.1400 1.7000 ;
        RECT 6.5650 1.3900 6.6550 1.6600 ;
    END
    ANTENNADIFFAREA 0.5616 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 6.2450 2.0350 6.4500 2.0800 ;
        RECT 5.2600 2.0300 5.4700 2.0800 ;
        RECT 3.9250 2.0250 4.1350 2.0800 ;
        RECT 5.7850 2.0200 5.8750 2.0800 ;
        RECT 1.0250 1.9850 1.1450 2.0800 ;
        RECT 7.0800 1.7300 7.2500 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 1.0450 1.5500 1.4150 ;
    END
    ANTENNAGATEAREA 0.0816 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9800 1.4650 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2400 0.8950 7.3500 1.3050 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 1.6800 0.4800 6.9050 0.5700 ;
      RECT 6.8150 0.5700 6.9050 1.4600 ;
      RECT 3.9500 0.5700 4.0400 1.0650 ;
      RECT 4.3900 0.5700 4.4800 1.5350 ;
      RECT 1.6600 1.2850 1.7700 1.4550 ;
      RECT 1.6800 0.5700 1.7700 1.2850 ;
      RECT 1.9250 0.4600 2.0950 0.4800 ;
      RECT 6.7600 1.5500 7.5300 1.6400 ;
      RECT 7.4100 1.4500 7.5300 1.5500 ;
      RECT 7.4400 0.7000 7.5300 1.4500 ;
      RECT 7.4100 0.5300 7.5300 0.7000 ;
      RECT 7.0150 1.0000 7.1050 1.5500 ;
      RECT 1.8650 1.8300 6.8500 1.9200 ;
      RECT 6.7600 1.6400 6.8500 1.8300 ;
      RECT 3.9500 1.3350 4.0400 1.8300 ;
      RECT 4.7500 0.8850 4.8400 1.8300 ;
      RECT 0.3350 1.8800 0.7500 1.9700 ;
      RECT 0.3350 1.7900 0.4250 1.8800 ;
      RECT 0.0600 1.7000 0.4250 1.7900 ;
      RECT 0.0600 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5200 0.5100 0.6000 ;
      RECT 0.4200 0.4300 0.8300 0.5200 ;
      RECT 0.0600 0.6900 0.1500 1.7000 ;
      RECT 0.5150 1.7000 1.6300 1.7900 ;
      RECT 0.4450 0.8100 1.5900 0.9000 ;
      RECT 1.5000 0.4900 1.5900 0.8100 ;
      RECT 1.0700 0.9000 1.1600 1.7000 ;
      RECT 0.5150 1.5450 0.6050 1.7000 ;
      RECT 0.4450 0.9000 0.6550 0.9350 ;
      RECT 1.7250 1.5900 1.9500 1.6800 ;
      RECT 1.8600 1.1500 1.9500 1.5900 ;
      RECT 1.8600 1.0600 2.8250 1.1500 ;
      RECT 2.7350 1.1500 2.8250 1.2950 ;
      RECT 1.8600 0.6800 1.9500 1.0600 ;
      RECT 2.6000 0.6700 3.3300 0.7600 ;
      RECT 2.1850 1.6400 3.5900 1.7300 ;
      RECT 3.5000 0.9400 3.5900 1.6400 ;
      RECT 2.8600 0.8500 3.5900 0.9400 ;
      RECT 2.1850 1.2550 2.2750 1.6400 ;
      RECT 4.5700 0.6700 5.4900 0.7600 ;
      RECT 5.4000 0.7600 5.4900 1.1350 ;
      RECT 4.1500 1.6450 4.6600 1.7350 ;
      RECT 4.1500 1.2450 4.2400 1.6450 ;
      RECT 4.5700 0.7600 4.6600 1.6450 ;
      RECT 3.7200 1.1550 4.2400 1.2450 ;
      RECT 3.7200 1.2450 3.8100 1.6300 ;
      RECT 3.7200 0.7750 3.8100 1.1550 ;
      RECT 5.5800 1.0650 6.3000 1.1550 ;
      RECT 4.9300 1.6500 5.6700 1.7400 ;
      RECT 5.5800 1.1550 5.6700 1.6500 ;
      RECT 5.5800 0.6800 5.6700 1.0650 ;
      RECT 4.9300 1.3700 5.0200 1.6500 ;
  END
END SDFFSRPQ_X3M_A12TH

MACRO SDFFSRPQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.0750 0.3200 0.2150 0.4650 ;
        RECT 1.0350 0.3200 1.1350 0.6500 ;
        RECT 4.3250 0.3200 4.4150 0.3600 ;
        RECT 5.5450 0.3200 5.7550 0.3900 ;
        RECT 6.0700 0.3200 6.2750 0.3900 ;
        RECT 6.5900 0.3200 6.7900 0.3700 ;
        RECT 7.1200 0.3200 7.4950 0.3450 ;
        RECT 7.6750 0.3200 7.8450 0.8250 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 1.0450 1.5500 1.4150 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9600 1.4650 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4100 1.4600 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 1.1000 4.3700 1.5000 ;
    END
    ANTENNAGATEAREA 0.135 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2100 1.0400 5.5450 1.1800 ;
    END
    ANTENNAGATEAREA 0.123 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.3450 0.8500 7.0350 0.9500 ;
        RECT 6.8500 0.9500 6.9500 1.3000 ;
        RECT 6.3450 0.7150 6.5150 0.8500 ;
        RECT 6.8650 0.7150 7.0350 0.8500 ;
        RECT 6.3800 1.3000 7.0000 1.4000 ;
        RECT 6.3800 1.4000 6.4800 1.7150 ;
        RECT 6.9000 1.4000 7.0000 1.7000 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 3.0950 2.0500 3.2850 2.0800 ;
        RECT 4.0950 2.0500 4.2650 2.0800 ;
        RECT 6.0850 2.0350 6.2950 2.0800 ;
        RECT 6.5850 2.0350 6.7900 2.0800 ;
        RECT 5.5450 2.0300 5.7550 2.0800 ;
        RECT 1.0250 2.0150 1.1450 2.0800 ;
        RECT 7.7250 1.7200 7.8350 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6950 1.0100 7.9500 1.1200 ;
        RECT 7.8500 1.1200 7.9500 1.3200 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 2.1650 1.6400 3.5450 1.7300 ;
      RECT 2.1650 1.2350 2.2550 1.6400 ;
      RECT 3.4550 0.9400 3.5450 1.6400 ;
      RECT 2.8550 0.8500 3.5450 0.9400 ;
      RECT 3.4550 0.7800 3.5450 0.8500 ;
      RECT 3.4550 0.6900 3.9300 0.7800 ;
      RECT 4.7850 0.6700 5.7350 0.7600 ;
      RECT 5.6450 0.7600 5.7350 0.9950 ;
      RECT 5.6450 0.9950 5.7950 1.1650 ;
      RECT 3.6450 1.6450 4.8750 1.7350 ;
      RECT 4.7850 0.7600 4.8750 1.6450 ;
      RECT 3.6450 1.0550 3.7350 1.6450 ;
      RECT 3.6450 0.9650 4.1500 1.0550 ;
      RECT 4.0600 0.7250 4.1500 0.9650 ;
      RECT 5.9650 1.0650 6.6400 1.1550 ;
      RECT 5.1650 1.6400 6.0550 1.7300 ;
      RECT 5.1650 1.3700 5.2550 1.6400 ;
      RECT 5.9650 1.1550 6.0550 1.6400 ;
      RECT 5.9650 0.7700 6.0550 1.0650 ;
      RECT 5.8250 0.6800 6.0550 0.7700 ;
      RECT 1.7000 0.4800 7.5200 0.5700 ;
      RECT 7.4300 0.5700 7.5200 1.4500 ;
      RECT 4.5850 0.5700 4.6750 1.5450 ;
      RECT 1.7000 0.5700 1.7900 1.4550 ;
      RECT 7.2300 1.5400 8.1300 1.6300 ;
      RECT 8.0150 1.4500 8.1300 1.5400 ;
      RECT 8.0400 0.8150 8.1300 1.4500 ;
      RECT 8.0150 0.4450 8.1300 0.8150 ;
      RECT 1.9200 1.8300 7.3200 1.9200 ;
      RECT 7.2300 1.6300 7.3200 1.8300 ;
      RECT 7.2300 1.1850 7.3200 1.5400 ;
      RECT 7.2300 1.0150 7.3350 1.1850 ;
      RECT 4.9850 0.8850 5.0750 1.8300 ;
      RECT 0.3350 1.8800 0.7500 1.9700 ;
      RECT 0.3350 1.7900 0.4250 1.8800 ;
      RECT 0.0600 1.7000 0.4250 1.7900 ;
      RECT 0.0600 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5200 0.5100 0.6000 ;
      RECT 0.4200 0.4300 0.8100 0.5200 ;
      RECT 0.0600 0.6900 0.1500 1.7000 ;
      RECT 1.4600 1.7900 1.6300 1.9900 ;
      RECT 0.5150 1.7000 1.6300 1.7900 ;
      RECT 0.4450 0.8450 1.5900 0.9350 ;
      RECT 1.5000 0.5250 1.5900 0.8450 ;
      RECT 1.0600 0.9350 1.1500 1.7000 ;
      RECT 0.5150 1.5450 0.6050 1.7000 ;
      RECT 1.7250 1.5900 1.9700 1.6800 ;
      RECT 1.8800 0.9600 1.9700 1.5900 ;
      RECT 1.8800 0.8700 2.7450 0.9600 ;
      RECT 2.6550 0.9600 2.7450 1.1000 ;
      RECT 1.8800 0.7000 1.9700 0.8700 ;
      RECT 2.6550 1.1000 2.8700 1.1900 ;
      RECT 2.5750 0.6700 3.3050 0.7600 ;
      RECT 2.4500 1.4350 3.3500 1.5250 ;
      RECT 2.4500 1.0600 2.5400 1.4350 ;
      RECT 3.2600 1.0550 3.3500 1.4350 ;
  END
END SDFFSRPQ_X4M_A12TH

MACRO SDFFYQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.9400 ;
        RECT 0.9900 0.3200 1.1600 0.6050 ;
        RECT 2.4100 0.3200 2.5800 0.5600 ;
        RECT 4.4350 0.3200 4.6050 0.3750 ;
        RECT 4.9650 0.3200 5.0650 0.7300 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8900 5.1500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9700 4.3500 1.2900 ;
        RECT 4.1550 1.2900 4.3500 1.3900 ;
        RECT 4.1650 0.8700 4.3500 0.9700 ;
        RECT 4.1550 1.3900 4.2550 1.7100 ;
        RECT 4.1650 0.7450 4.2650 0.8700 ;
    END
    ANTENNADIFFAREA 0.26455 ;
  END Q

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.2500 0.8700 1.3500 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 3.4150 2.0250 3.6250 2.0800 ;
        RECT 2.2800 1.9900 2.4500 2.0800 ;
        RECT 1.0700 1.8800 1.1800 2.0800 ;
        RECT 0.3350 1.6650 0.4450 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0500 1.3700 1.4200 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 1.4500 0.7900 1.5700 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI
  OBS
    LAYER M1 ;
      RECT 0.0450 1.0350 1.1350 1.1250 ;
      RECT 0.9300 1.1250 1.1350 1.1550 ;
      RECT 0.0450 1.6550 0.1950 1.8400 ;
      RECT 0.0450 1.1250 0.1350 1.6550 ;
      RECT 0.0850 0.8100 0.1750 1.0350 ;
      RECT 0.7700 1.7000 1.6700 1.7900 ;
      RECT 1.5000 0.9400 1.5900 1.7000 ;
      RECT 0.7850 0.8500 1.5900 0.9400 ;
      RECT 1.5000 0.6150 1.5900 0.8500 ;
      RECT 1.7600 1.6100 1.9750 1.7000 ;
      RECT 1.8850 1.4450 1.9750 1.6100 ;
      RECT 1.8850 1.3550 2.5300 1.4450 ;
      RECT 1.8850 0.6800 1.9750 1.3550 ;
      RECT 2.6300 1.1850 2.7200 1.6150 ;
      RECT 2.2000 1.0950 2.8100 1.1850 ;
      RECT 2.7200 0.9500 2.8100 1.0950 ;
      RECT 2.7200 0.8600 2.9600 0.9500 ;
      RECT 2.8800 1.6200 3.1600 1.7100 ;
      RECT 3.0700 0.7850 3.1600 1.6200 ;
      RECT 3.0700 0.6950 3.5200 0.7850 ;
      RECT 3.4300 0.7850 3.5200 1.1300 ;
      RECT 3.4300 1.1300 3.8150 1.2400 ;
      RECT 3.9650 1.0850 4.1600 1.1750 ;
      RECT 3.7050 1.6200 4.0550 1.7100 ;
      RECT 3.9650 1.4350 4.0550 1.6200 ;
      RECT 3.4300 1.3450 4.0550 1.4350 ;
      RECT 3.4300 1.4350 3.5200 1.5350 ;
      RECT 3.9650 1.1750 4.0550 1.3450 ;
      RECT 3.9650 0.7700 4.0550 1.0850 ;
      RECT 3.8600 0.6800 4.0550 0.7700 ;
      RECT 4.4400 1.6500 4.8700 1.7400 ;
      RECT 4.4400 0.9000 4.5300 1.6500 ;
      RECT 4.4400 0.8100 4.8900 0.9000 ;
      RECT 4.4400 0.5700 4.5300 0.8100 ;
      RECT 2.7400 0.4800 4.5300 0.5700 ;
      RECT 2.7400 0.5700 2.8300 0.6800 ;
      RECT 2.1250 0.6800 2.8300 0.7700 ;
      RECT 2.1250 0.5700 2.2150 0.6800 ;
      RECT 1.6850 0.4800 2.2150 0.5700 ;
      RECT 1.6850 0.5700 1.7750 1.5000 ;
      RECT 2.5750 1.9000 5.3300 1.9200 ;
      RECT 1.9000 1.8300 5.3300 1.9000 ;
      RECT 5.2300 1.5600 5.3300 1.8300 ;
      RECT 4.6250 1.4700 5.3300 1.5600 ;
      RECT 5.2400 0.7800 5.3300 1.4700 ;
      RECT 5.1900 0.5700 5.3300 0.7800 ;
      RECT 4.6250 1.0150 4.7150 1.4700 ;
      RECT 1.9000 1.8100 2.6650 1.8300 ;
      RECT 3.2500 1.0100 3.3400 1.8300 ;
  END
END SDFFYQ_X1M_A12TH

MACRO SDFFYQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.9400 ;
        RECT 0.9900 0.3200 1.1600 0.6050 ;
        RECT 2.4550 0.3200 2.6250 0.5600 ;
        RECT 3.5900 0.3200 3.7600 0.3800 ;
        RECT 4.1650 0.3200 4.3350 0.3700 ;
        RECT 4.6850 0.3200 4.8550 0.3700 ;
        RECT 5.6000 0.3200 5.7000 0.8050 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 1.4500 0.7900 1.5700 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 0.9150 5.5600 1.3500 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.2500 0.8700 1.3500 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7250 4.5600 1.7050 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 2.2150 1.9900 2.3850 2.0800 ;
        RECT 1.0700 1.8800 1.1800 2.0800 ;
        RECT 0.3350 1.6650 0.4450 2.0800 ;
        RECT 5.6300 1.5000 5.7200 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0500 1.3700 1.4200 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.0450 1.0350 1.1350 1.1250 ;
      RECT 0.9300 1.1250 1.1350 1.1550 ;
      RECT 0.0450 1.6550 0.1950 1.8400 ;
      RECT 0.0450 1.1250 0.1350 1.6550 ;
      RECT 0.0850 0.7900 0.1750 1.0350 ;
      RECT 0.7700 1.7000 1.6700 1.7900 ;
      RECT 1.5000 0.9400 1.5900 1.7000 ;
      RECT 0.7850 0.8500 1.5900 0.9400 ;
      RECT 1.5000 0.6150 1.5900 0.8500 ;
      RECT 1.7600 1.5850 1.9750 1.6750 ;
      RECT 1.8850 1.3700 1.9750 1.5850 ;
      RECT 1.8850 1.2800 2.4700 1.3700 ;
      RECT 2.3800 1.3700 2.4700 1.4800 ;
      RECT 1.8850 0.6800 1.9750 1.2800 ;
      RECT 2.5800 1.1600 2.6700 1.7050 ;
      RECT 2.2000 1.0700 2.8100 1.1600 ;
      RECT 2.7200 0.9500 2.8100 1.0700 ;
      RECT 2.7200 0.8600 2.9850 0.9500 ;
      RECT 2.9650 1.3000 3.0550 1.7400 ;
      RECT 2.9650 1.2100 3.2100 1.3000 ;
      RECT 3.1200 0.8800 3.2100 1.2100 ;
      RECT 3.1200 0.7900 3.6300 0.8800 ;
      RECT 3.5400 0.8800 3.6300 0.9850 ;
      RECT 3.5400 0.9850 3.8700 1.0750 ;
      RECT 3.7800 1.0750 3.8700 1.2300 ;
      RECT 3.8250 1.6200 4.0800 1.7100 ;
      RECT 3.9900 1.4350 4.0800 1.6200 ;
      RECT 3.4800 1.3450 4.0800 1.4350 ;
      RECT 3.4800 1.4350 3.5700 1.5350 ;
      RECT 3.9900 1.1950 4.0800 1.3450 ;
      RECT 3.9900 1.0250 4.1600 1.1950 ;
      RECT 3.9900 0.8300 4.0900 1.0250 ;
      RECT 3.8950 0.7300 4.0900 0.8300 ;
      RECT 5.0350 1.3600 5.1250 1.7000 ;
      RECT 4.7150 1.2700 5.1250 1.3600 ;
      RECT 4.7150 0.5700 4.8050 1.2700 ;
      RECT 2.7400 0.4800 5.1800 0.5700 ;
      RECT 5.0900 0.5700 5.1800 0.9350 ;
      RECT 2.7400 0.5700 2.8300 0.6800 ;
      RECT 3.2100 0.4100 3.3800 0.4800 ;
      RECT 2.1250 0.6800 2.8300 0.7700 ;
      RECT 2.1250 0.5700 2.2150 0.6800 ;
      RECT 1.6850 0.4800 2.2150 0.5700 ;
      RECT 1.6850 0.5700 1.7750 1.4750 ;
      RECT 2.4500 1.9000 5.4350 1.9200 ;
      RECT 1.9000 1.8300 5.4350 1.9000 ;
      RECT 5.2700 1.5300 5.4350 1.8300 ;
      RECT 5.2700 1.1500 5.3600 1.5300 ;
      RECT 4.9150 1.0600 5.3600 1.1500 ;
      RECT 5.2700 0.8050 5.3600 1.0600 ;
      RECT 5.2700 0.7150 5.4350 0.8050 ;
      RECT 5.3450 0.4200 5.4350 0.7150 ;
      RECT 1.9000 1.8100 2.5400 1.8300 ;
      RECT 2.7600 1.3150 2.8500 1.8300 ;
      RECT 3.3000 1.0500 3.3900 1.8300 ;
  END
END SDFFYQ_X2M_A12TH

MACRO SDFFYQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0500 0.3200 0.2400 0.3500 ;
        RECT 0.9150 0.3200 1.0150 0.6100 ;
        RECT 1.9550 0.3200 2.3250 0.3750 ;
        RECT 3.3650 0.3200 3.5350 0.3600 ;
        RECT 3.9400 0.3200 4.1100 0.3750 ;
        RECT 4.4600 0.3200 4.6300 0.3600 ;
        RECT 5.3100 0.3200 5.4100 0.7300 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1950 0.9500 1.3900 ;
        RECT 0.7700 1.0100 0.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.9700 4.7500 1.3000 ;
        RECT 4.2350 1.3000 4.8550 1.4000 ;
        RECT 4.2000 0.8700 4.8550 0.9700 ;
        RECT 4.2350 1.4000 4.3350 1.7100 ;
        RECT 4.7550 1.4000 4.8550 1.7100 ;
        RECT 4.7550 0.7300 4.8550 0.8700 ;
        RECT 4.2000 0.6650 4.3700 0.8700 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4450 1.0200 5.5650 1.5000 ;
    END
    ANTENNAGATEAREA 0.0537 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0500 1.3600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0873 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0150 0.3600 1.4500 ;
    END
    ANTENNAGATEAREA 0.0747 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 1.9650 2.0100 2.3350 2.0800 ;
        RECT 0.8750 1.8350 1.0450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3950 0.4400 0.8000 0.5400 ;
      RECT 0.0500 1.8200 0.7500 1.9200 ;
      RECT 0.0500 0.5850 0.4950 0.6850 ;
      RECT 0.3950 0.5400 0.4950 0.5850 ;
      RECT 0.0500 0.6850 0.1500 1.8200 ;
      RECT 1.3350 1.7300 1.5050 1.9650 ;
      RECT 0.4500 1.6400 1.5050 1.7300 ;
      RECT 0.3800 0.8000 1.4700 0.9000 ;
      RECT 1.3700 0.4800 1.4700 0.8000 ;
      RECT 0.4500 0.9250 0.5400 1.6400 ;
      RECT 0.3800 0.9000 0.6950 0.9250 ;
      RECT 1.6450 1.5700 1.9100 1.6600 ;
      RECT 1.8200 1.0500 1.9100 1.5700 ;
      RECT 1.8200 0.9600 2.4500 1.0500 ;
      RECT 2.3600 1.0500 2.4500 1.2400 ;
      RECT 1.8200 0.8550 1.9100 0.9600 ;
      RECT 1.7400 0.6850 1.9100 0.8550 ;
      RECT 2.0650 1.5850 2.6300 1.6750 ;
      RECT 2.0650 1.1400 2.1550 1.5850 ;
      RECT 2.5400 0.7300 2.6300 1.5850 ;
      RECT 2.7250 0.9250 2.8150 1.7150 ;
      RECT 2.7250 0.8350 3.6150 0.9250 ;
      RECT 3.5250 0.9250 3.6150 1.2450 ;
      RECT 3.7300 1.0800 4.5350 1.1800 ;
      RECT 3.7300 1.4450 3.8200 1.7300 ;
      RECT 3.2900 1.3550 3.8200 1.4450 ;
      RECT 3.2900 1.2300 3.3800 1.3550 ;
      RECT 3.7300 1.1800 3.8200 1.3550 ;
      RECT 3.7300 0.7500 3.8200 1.0800 ;
      RECT 1.5600 0.4850 5.1000 0.5750 ;
      RECT 5.0100 0.5750 5.1000 1.6450 ;
      RECT 1.5600 1.3250 1.7300 1.4350 ;
      RECT 1.5600 0.5750 1.6500 1.3250 ;
      RECT 3.0550 0.4400 3.2250 0.4850 ;
      RECT 1.7500 1.8300 5.7550 1.9200 ;
      RECT 5.5850 1.6300 5.7550 1.8300 ;
      RECT 5.6650 0.9300 5.7550 1.6300 ;
      RECT 5.1950 0.8400 5.7550 0.9300 ;
      RECT 5.6250 0.5200 5.7550 0.8400 ;
      RECT 5.1950 0.9300 5.2850 1.2600 ;
      RECT 3.0600 1.0250 3.1500 1.8300 ;
  END
END SDFFYQ_X3M_A12TH

MACRO RF2R1WS_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.9150 ;
        RECT 0.6400 0.3200 0.7400 0.5600 ;
        RECT 2.3800 0.3200 2.7500 0.3750 ;
        RECT 3.1900 0.3200 3.2900 0.5050 ;
        RECT 4.4700 0.3200 4.6800 0.3850 ;
        RECT 5.5650 0.3200 5.6650 0.6550 ;
    END
  END VSS

  PIN WWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.2500 1.1500 ;
    END
    ANTENNAGATEAREA 0.1146 ;
  END WWL

  PIN RBL2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9550 1.0500 5.3150 1.1500 ;
        RECT 4.9550 1.1500 5.0550 1.5600 ;
        RECT 4.9550 0.7600 5.0550 1.0500 ;
        RECT 4.9550 1.5600 5.2000 1.6600 ;
        RECT 4.9550 0.6600 5.1900 0.7600 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END RBL2

  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 1.1450 3.7500 1.4900 ;
        RECT 3.6500 1.4900 3.7750 1.7100 ;
        RECT 3.6500 1.0450 3.8000 1.1450 ;
        RECT 3.7000 0.8100 3.8000 1.0450 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END RBL1

  PIN RWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1650 0.8500 5.7600 0.9500 ;
        RECT 5.6600 0.9500 5.7600 1.2400 ;
    END
    ANTENNAGATEAREA 0.1044 ;
  END RWL2

  PIN RWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3650 1.2100 4.5500 1.3800 ;
        RECT 4.4500 1.3800 4.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.1044 ;
  END RWL1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 0.6100 1.8400 0.7100 2.0800 ;
        RECT 0.0900 1.7750 0.1900 2.0800 ;
        RECT 4.5250 1.7050 4.6250 2.0800 ;
        RECT 5.5650 1.7050 5.6650 2.0800 ;
        RECT 3.1600 1.4950 3.2600 2.0800 ;
    END
  END VDD

  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1400 0.1600 1.6000 ;
    END
    ANTENNAGATEAREA 0.1308 ;
  END WBL
  OBS
    LAYER M1 ;
      RECT 0.3550 1.6500 1.6500 1.7400 ;
      RECT 0.3550 0.6700 1.6500 0.7600 ;
      RECT 0.3550 1.7400 0.4450 1.9700 ;
      RECT 0.3550 0.7600 0.4450 1.6500 ;
      RECT 0.9750 1.3400 1.0650 1.5000 ;
      RECT 0.9750 1.2500 1.7950 1.3400 ;
      RECT 1.7050 0.9400 1.7950 1.2500 ;
      RECT 0.9000 0.8500 2.1200 0.9400 ;
      RECT 1.9250 0.8000 2.1200 0.8500 ;
      RECT 2.3550 1.1750 2.4450 1.4700 ;
      RECT 2.1600 1.0850 2.4450 1.1750 ;
      RECT 2.3550 0.8050 2.4450 1.0850 ;
      RECT 3.4200 1.8200 4.0500 1.9100 ;
      RECT 3.9600 1.6200 4.0500 1.8200 ;
      RECT 3.9600 1.5200 4.0550 1.6200 ;
      RECT 3.9650 0.7850 4.0550 1.5200 ;
      RECT 3.4200 1.3450 3.5100 1.8200 ;
      RECT 2.9050 1.2550 3.5100 1.3450 ;
      RECT 3.4200 0.9750 3.5100 1.2550 ;
      RECT 3.4200 0.8050 3.5350 0.9750 ;
      RECT 2.9050 1.3450 2.9950 1.7200 ;
      RECT 2.9050 0.7950 2.9950 1.2550 ;
      RECT 4.2100 1.6100 4.3000 1.9300 ;
      RECT 4.1450 1.5200 4.3000 1.6100 ;
      RECT 4.1450 0.8300 4.2350 1.5200 ;
      RECT 4.1450 0.7400 4.3600 0.8300 ;
      RECT 3.6100 0.5050 4.6450 0.5950 ;
      RECT 4.5550 0.5950 4.6450 1.1000 ;
      RECT 2.1750 0.6050 3.7000 0.6950 ;
      RECT 3.6100 0.5950 3.7000 0.6050 ;
      RECT 2.0550 1.5800 2.7200 1.6700 ;
      RECT 2.0550 1.5600 2.1450 1.5800 ;
      RECT 2.6300 0.6950 2.7200 1.5800 ;
      RECT 1.1800 1.4700 2.1450 1.5600 ;
      RECT 2.1750 0.5700 2.2650 0.6050 ;
      RECT 1.1800 0.4800 2.2650 0.5700 ;
      RECT 4.7350 1.8300 5.4000 1.9200 ;
      RECT 5.3100 1.5300 5.4000 1.8300 ;
      RECT 4.7350 0.4800 5.4600 0.5700 ;
      RECT 4.7350 0.5700 4.8250 1.8300 ;
      RECT 5.8300 1.4400 5.9200 1.9050 ;
      RECT 5.2050 1.3500 5.9550 1.4400 ;
      RECT 5.8650 0.7450 5.9550 1.3500 ;
      RECT 5.8100 0.5750 5.9550 0.7450 ;
      RECT 5.2050 1.2550 5.2950 1.3500 ;
  END
END RF2R1WS_X1P4M_A12TH

MACRO RF2R1WS_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7500 ;
        RECT 0.6050 0.3200 0.7750 0.5800 ;
        RECT 2.3800 0.3200 2.7500 0.3750 ;
        RECT 3.1600 0.3200 3.2600 0.4350 ;
        RECT 4.9900 0.3200 5.0900 0.6650 ;
    END
  END VSS

  PIN RBL2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.8950 5.9500 1.5850 ;
        RECT 5.7050 1.5850 5.9500 1.6750 ;
        RECT 5.7050 0.7950 5.9500 0.8950 ;
    END
    ANTENNADIFFAREA 0.286 ;
  END RBL2

  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.7600 3.7650 1.7100 ;
    END
    ANTENNADIFFAREA 0.286 ;
  END RBL1

  PIN RWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2400 1.0500 5.7100 1.1500 ;
    END
    ANTENNAGATEAREA 0.1452 ;
  END RWL2

  PIN RWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3600 1.2100 4.5500 1.3100 ;
        RECT 4.4500 1.3100 4.5500 1.5550 ;
        RECT 4.3600 1.0000 4.4600 1.2100 ;
    END
    ANTENNAGATEAREA 0.1452 ;
  END RWL1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.6100 1.8300 0.7100 2.0800 ;
        RECT 0.0900 1.7900 0.1900 2.0800 ;
        RECT 3.1600 1.7700 3.2600 2.0800 ;
        RECT 4.4700 1.7700 4.5700 2.0800 ;
        RECT 4.9550 1.7200 5.1250 2.0800 ;
    END
  END VDD

  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2400 0.1500 1.6000 ;
        RECT 0.0500 1.0700 0.2650 1.2400 ;
    END
    ANTENNAGATEAREA 0.1872 ;
  END WBL

  PIN WWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8450 1.0500 1.2650 1.1700 ;
    END
    ANTENNAGATEAREA 0.1518 ;
  END WWL
  OBS
    LAYER M1 ;
      RECT 1.4600 1.7400 1.6300 1.9600 ;
      RECT 0.3550 1.6500 1.6300 1.7400 ;
      RECT 0.3550 0.6700 1.6500 0.7600 ;
      RECT 0.3550 0.7600 0.4450 1.6500 ;
      RECT 0.3550 0.5400 0.4450 0.6700 ;
      RECT 0.9750 1.3500 1.0650 1.5000 ;
      RECT 0.9750 1.2600 1.7950 1.3500 ;
      RECT 1.7050 0.9400 1.7950 1.2600 ;
      RECT 0.9150 0.8500 2.1200 0.9400 ;
      RECT 1.9250 0.8000 2.1200 0.8500 ;
      RECT 2.3550 1.1750 2.4450 1.4700 ;
      RECT 2.1600 1.0850 2.4450 1.1750 ;
      RECT 2.3550 0.8050 2.4450 1.0850 ;
      RECT 3.4150 1.8200 4.0250 1.9100 ;
      RECT 3.9350 0.7600 4.0250 1.8200 ;
      RECT 3.4150 1.3450 3.5050 1.8200 ;
      RECT 2.9050 1.2550 3.5050 1.3450 ;
      RECT 3.4150 0.7850 3.5050 1.2550 ;
      RECT 2.9050 1.3450 2.9950 1.7200 ;
      RECT 2.9050 0.7850 2.9950 1.2550 ;
      RECT 4.1400 1.6700 4.3350 1.9600 ;
      RECT 4.1400 0.7500 4.2300 1.6700 ;
      RECT 4.1400 0.6600 4.3350 0.7500 ;
      RECT 3.3750 0.4800 4.6400 0.5700 ;
      RECT 4.5500 0.5700 4.6400 1.0250 ;
      RECT 4.5500 1.0250 4.7900 1.1150 ;
      RECT 1.7600 1.6700 1.8500 1.9000 ;
      RECT 1.7600 1.5800 2.7200 1.6700 ;
      RECT 1.7600 1.5600 1.8500 1.5800 ;
      RECT 2.6300 0.6850 2.7200 1.5800 ;
      RECT 1.1900 1.4700 1.8500 1.5600 ;
      RECT 2.1750 0.5700 2.2650 0.5950 ;
      RECT 1.1800 0.4800 2.2650 0.5700 ;
      RECT 2.1750 0.5950 3.4650 0.6850 ;
      RECT 3.3750 0.5700 3.4650 0.5950 ;
      RECT 5.0600 1.3500 5.6450 1.4400 ;
      RECT 5.5550 1.2500 5.6450 1.3500 ;
      RECT 5.0600 0.7950 5.3450 0.8850 ;
      RECT 5.2550 0.4950 5.3450 0.7950 ;
      RECT 5.0600 0.8850 5.1500 1.3500 ;
      RECT 5.5050 1.7650 6.1300 1.8550 ;
      RECT 6.0250 1.8550 6.1300 1.9550 ;
      RECT 6.0400 0.6450 6.1300 1.7650 ;
      RECT 5.5050 0.5550 6.1300 0.6450 ;
      RECT 6.0250 0.4150 6.1300 0.5550 ;
      RECT 5.5050 1.8550 5.5950 1.9750 ;
      RECT 5.5050 1.6200 5.5950 1.7650 ;
      RECT 4.7350 1.5300 5.5950 1.6200 ;
      RECT 5.5050 0.6450 5.5950 0.8350 ;
      RECT 5.5050 0.4100 5.5950 0.5550 ;
      RECT 4.8800 0.8950 4.9700 1.5300 ;
      RECT 4.7350 0.8050 4.9700 0.8950 ;
      RECT 4.7350 1.6200 4.8250 1.9600 ;
      RECT 4.7350 0.4850 4.8250 0.8050 ;
  END
END RF2R1WS_X2M_A12TH

MACRO RF2R2WS_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 2.4800 0.3200 2.5700 0.3900 ;
        RECT 3.6700 0.3200 3.8400 0.3750 ;
        RECT 4.7900 0.3200 4.8900 0.9700 ;
        RECT 5.8300 0.3200 5.9200 0.6450 ;
    END
  END VSS

  PIN WBL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0050 0.5550 1.4300 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END WBL1

  PIN WWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.7500 3.5500 1.0750 ;
        RECT 3.3050 1.0750 3.5500 1.1650 ;
        RECT 1.7850 0.6600 3.5500 0.7500 ;
        RECT 1.7850 0.7500 1.8750 1.4650 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END WWL2

  PIN WBL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0050 2.7500 1.5450 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END WBL2

  PIN RBL2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9500 4.3500 1.5300 ;
        RECT 4.2500 1.5300 4.3650 1.7000 ;
        RECT 4.2500 0.5800 4.3650 0.9500 ;
    END
    ANTENNADIFFAREA 0.2288 ;
  END RBL2

  PIN WWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8950 0.3500 1.2250 ;
        RECT 0.2350 0.8050 0.5450 0.8950 ;
        RECT 0.4550 0.5700 0.5450 0.8050 ;
        RECT 0.4550 0.4800 0.9400 0.5700 ;
        RECT 0.8500 0.5700 0.9400 0.9200 ;
        RECT 0.8500 0.9200 1.2000 1.0100 ;
        RECT 1.1100 1.0100 1.2000 1.6900 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END WWL1

  PIN RWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6400 1.0550 4.7500 1.4700 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END RWL2

  PIN RWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.3800 4.9500 1.6200 ;
        RECT 4.8500 1.2100 4.9850 1.3800 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END RWL1

  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2100 0.6100 5.4100 0.7500 ;
        RECT 5.3100 0.7500 5.4100 1.7200 ;
    END
    ANTENNADIFFAREA 0.2288 ;
  END RBL1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6700 0.6900 0.7600 1.4700 ;
      RECT 0.0550 1.6450 0.9400 1.7350 ;
      RECT 0.8500 1.2400 0.9400 1.6450 ;
      RECT 0.8500 1.1500 1.0200 1.2400 ;
      RECT 0.0550 1.4850 0.1700 1.6450 ;
      RECT 0.0550 0.7400 0.1450 1.4850 ;
      RECT 0.0550 0.5700 0.1700 0.7400 ;
      RECT 1.5550 1.5900 2.4600 1.6800 ;
      RECT 2.2250 0.9550 2.3150 1.5900 ;
      RECT 2.2250 0.8650 2.4800 0.9550 ;
      RECT 1.5550 1.0100 1.6450 1.5900 ;
      RECT 2.8650 1.2900 2.9950 1.4600 ;
      RECT 2.9050 0.9550 2.9950 1.2900 ;
      RECT 2.8250 0.8650 2.9950 0.9550 ;
      RECT 3.4050 1.4250 3.4950 1.7200 ;
      RECT 3.2650 1.3350 3.7400 1.4250 ;
      RECT 3.6500 0.5700 3.7400 1.3350 ;
      RECT 1.4700 0.4800 3.7400 0.5700 ;
      RECT 1.4700 0.5700 1.5600 0.8900 ;
      RECT 4.0100 0.5600 4.1200 1.6550 ;
      RECT 4.4600 1.6050 4.6650 1.6950 ;
      RECT 4.4600 0.8400 4.6550 0.9300 ;
      RECT 4.4600 1.4950 4.5500 1.6050 ;
      RECT 4.4550 1.3250 4.5500 1.4950 ;
      RECT 4.4600 0.9300 4.5500 1.3250 ;
      RECT 5.0600 1.5200 5.1500 1.7350 ;
      RECT 5.0600 1.4300 5.2200 1.5200 ;
      RECT 5.1300 0.9300 5.2200 1.4300 ;
      RECT 5.0200 0.8400 5.2200 0.9300 ;
      RECT 5.5700 0.6100 5.6600 1.6550 ;
      RECT 0.8900 1.8300 5.8450 1.9200 ;
      RECT 5.7550 1.9200 5.8450 1.9250 ;
      RECT 5.7550 1.0400 5.8450 1.8300 ;
      RECT 3.8300 1.0150 3.9200 1.8300 ;
      RECT 1.2900 0.8100 1.3800 1.8300 ;
      RECT 1.0350 0.7200 1.3800 0.8100 ;
      RECT 1.0350 0.4700 1.1250 0.7200 ;
      RECT 3.0850 1.5400 3.2450 1.8300 ;
      RECT 3.0850 0.9550 3.1750 1.5400 ;
      RECT 3.0850 0.8650 3.2850 0.9550 ;
      RECT 2.1400 1.9200 2.3100 1.9250 ;
  END
END RF2R2WS_X1M_A12TH

MACRO RF2R2WS_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.6450 0.3200 ;
        RECT 1.1300 0.3200 1.2200 0.6100 ;
        RECT 1.6550 0.3200 1.7450 0.6550 ;
        RECT 2.1750 0.3200 2.2650 0.4350 ;
        RECT 3.3550 0.3200 3.4450 0.3900 ;
        RECT 4.4250 0.3200 4.5950 0.5950 ;
        RECT 4.8700 0.3200 5.0750 0.5950 ;
        RECT 6.0950 0.3200 6.2900 0.3900 ;
        RECT 6.8400 0.3200 6.9300 0.7100 ;
        RECT 7.3600 0.3200 7.4500 0.5150 ;
    END
  END VSS

  PIN RWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0050 1.0250 1.2800 1.1950 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END RWL1

  PIN RWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.3100 0.8500 7.6450 0.9500 ;
        RECT 7.5550 0.9500 7.6450 1.0450 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END RWL2

  PIN WWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2450 1.0500 5.7300 1.1600 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END WWL2

  PIN WBL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8000 1.0300 2.2150 1.1550 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END WBL1

  PIN WBL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0350 1.2500 6.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END WBL2

  PIN WWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.5700 3.9500 1.5600 ;
        RECT 3.2950 0.4800 3.9500 0.5700 ;
        RECT 3.2950 0.5700 3.3850 1.2700 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END WWL1

  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.4300 1.1000 ;
        RECT 0.2500 1.1000 0.3500 1.3700 ;
        RECT 0.3300 0.6200 0.4300 1.0100 ;
        RECT 0.2500 1.3700 0.4300 1.4600 ;
        RECT 0.3300 1.4600 0.4300 1.6800 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END RBL1

  PIN RBL2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.4500 0.8900 8.5500 1.4300 ;
        RECT 8.4300 0.5700 8.5500 0.8900 ;
        RECT 8.4300 1.4300 8.5500 1.8350 ;
        RECT 7.9700 0.5150 8.5500 0.5700 ;
        RECT 7.9700 0.5700 8.0600 1.5700 ;
        RECT 7.8500 0.4800 8.5500 0.5150 ;
        RECT 7.8600 1.5700 8.0600 1.6700 ;
        RECT 7.8500 0.4100 8.0600 0.4800 ;
    END
    ANTENNADIFFAREA 0.304925 ;
  END RBL2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.6450 2.7200 ;
        RECT 2.2100 2.0250 2.4200 2.0800 ;
        RECT 7.3600 2.0100 7.4500 2.0800 ;
        RECT 6.2000 1.9750 6.2900 2.0800 ;
        RECT 1.0400 1.9700 1.2800 2.0800 ;
        RECT 4.7450 1.8850 4.9500 2.0800 ;
        RECT 4.3600 1.8600 4.5300 2.0800 ;
        RECT 6.8400 1.7300 6.9300 2.0800 ;
        RECT 1.6500 1.6700 1.7400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8250 1.4350 0.9150 1.6600 ;
      RECT 0.7200 1.2250 0.9150 1.4350 ;
      RECT 0.8250 0.7400 0.9150 1.2250 ;
      RECT 0.8250 0.5300 0.9400 0.7400 ;
      RECT 0.0700 1.7900 1.4800 1.8800 ;
      RECT 1.3900 0.5000 1.4800 1.7900 ;
      RECT 0.5400 0.9750 0.6300 1.7900 ;
      RECT 0.5400 0.8850 0.6900 0.9750 ;
      RECT 0.6000 0.6050 0.6900 0.8850 ;
      RECT 0.0700 1.5050 0.1700 1.7900 ;
      RECT 0.0700 0.9650 0.1600 1.5050 ;
      RECT 0.0700 0.5950 0.1700 0.9650 ;
      RECT 2.9050 1.6000 3.1500 1.6900 ;
      RECT 2.9050 0.6100 2.9950 1.6000 ;
      RECT 2.3850 0.5200 2.9950 0.6100 ;
      RECT 2.3850 0.6100 2.4750 0.6450 ;
      RECT 1.9150 0.6450 2.4750 0.7350 ;
      RECT 2.3850 0.7350 2.4750 1.4100 ;
      RECT 1.9150 0.4650 2.0050 0.6450 ;
      RECT 2.0100 1.4100 2.5900 1.5000 ;
      RECT 2.0100 1.5000 2.1000 1.6650 ;
      RECT 2.5000 1.5000 2.5900 1.7400 ;
      RECT 3.2450 1.6500 3.4350 1.7400 ;
      RECT 3.2450 1.4700 3.3350 1.6500 ;
      RECT 3.0950 1.3800 3.5650 1.4700 ;
      RECT 3.4750 0.8600 3.5650 1.3800 ;
      RECT 3.0950 0.4300 3.1850 1.3800 ;
      RECT 4.4900 0.9550 4.5800 1.5900 ;
      RECT 4.2900 0.8650 4.7500 0.9550 ;
      RECT 5.0550 1.3100 5.7250 1.4000 ;
      RECT 5.0550 0.7850 5.3600 0.8750 ;
      RECT 5.0550 1.4000 5.1500 1.5900 ;
      RECT 5.0550 0.8750 5.1500 1.3100 ;
      RECT 5.0550 0.7750 5.1500 0.7850 ;
      RECT 4.0600 0.6850 5.1500 0.7750 ;
      RECT 4.0600 0.7750 4.1500 1.0550 ;
      RECT 5.2850 1.5850 6.5500 1.6750 ;
      RECT 6.4600 1.4750 6.5500 1.5850 ;
      RECT 5.4500 0.8700 6.5500 0.9600 ;
      RECT 5.9700 0.6800 6.0600 0.8700 ;
      RECT 6.4600 0.6600 6.5500 0.8700 ;
      RECT 5.8350 0.9600 5.9250 1.5850 ;
      RECT 5.4500 0.4100 5.5400 0.8700 ;
      RECT 6.6600 1.3150 7.3000 1.4050 ;
      RECT 1.8300 1.4450 1.9200 1.8300 ;
      RECT 1.5700 1.3550 1.9200 1.4450 ;
      RECT 1.5700 1.1850 1.6600 1.3550 ;
      RECT 2.7000 1.0150 2.7900 1.8300 ;
      RECT 2.6450 0.9250 2.7900 1.0150 ;
      RECT 2.6450 0.7450 2.7350 0.9250 ;
      RECT 3.7500 1.9200 3.8400 1.9850 ;
      RECT 1.8300 1.8300 3.8400 1.9200 ;
      RECT 3.6700 1.7700 3.8400 1.8300 ;
      RECT 3.6700 0.7500 3.7600 1.6800 ;
      RECT 3.5700 0.6600 3.7600 0.7500 ;
      RECT 4.7050 1.1300 4.7950 1.6800 ;
      RECT 5.7100 0.5700 5.8000 0.7800 ;
      RECT 5.7100 0.4100 5.8000 0.4800 ;
      RECT 3.6700 1.6800 5.1500 1.7700 ;
      RECT 5.0600 1.7700 5.1500 1.7950 ;
      RECT 5.0600 1.7950 6.7500 1.8850 ;
      RECT 6.6600 1.4050 6.7500 1.7950 ;
      RECT 6.6600 0.5700 6.7500 1.3150 ;
      RECT 5.7100 0.4800 6.7500 0.5700 ;
      RECT 7.6600 1.3250 7.8800 1.4150 ;
      RECT 7.7900 0.7600 7.8800 1.3250 ;
      RECT 7.6500 0.6700 7.8800 0.7600 ;
      RECT 7.6600 1.4150 7.7500 1.7400 ;
      RECT 7.4100 1.8300 8.2600 1.9200 ;
      RECT 8.1700 0.6600 8.2600 1.8300 ;
      RECT 7.1000 1.5200 7.5000 1.6100 ;
      RECT 7.4100 1.6100 7.5000 1.8300 ;
      RECT 7.4100 1.2250 7.5000 1.5200 ;
      RECT 7.1000 1.1350 7.5000 1.2250 ;
      RECT 7.1000 1.6100 7.1900 1.9700 ;
      RECT 7.1000 0.4100 7.1900 1.1350 ;
  END
END RF2R2WS_X1P4M_A12TH

MACRO RF2R2WS_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.6450 0.3200 ;
        RECT 1.1900 0.3200 1.2800 0.5800 ;
        RECT 1.7250 0.3200 1.8150 0.5800 ;
        RECT 2.2450 0.3200 2.3350 0.5800 ;
        RECT 3.4800 0.3200 3.5700 0.5950 ;
        RECT 4.2950 0.3200 4.4900 0.4150 ;
        RECT 4.8650 0.3200 5.0700 0.4100 ;
        RECT 6.2000 0.3200 6.2900 0.3900 ;
        RECT 6.8400 0.3200 6.9300 0.5600 ;
        RECT 7.3950 0.3200 7.4850 0.8550 ;
    END
  END VSS

  PIN RWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9750 1.1500 1.5950 ;
    END
    ANTENNAGATEAREA 0.144 ;
  END RWL1

  PIN RWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.9850 7.5700 1.4150 ;
    END
    ANTENNAGATEAREA 0.144 ;
  END RWL2

  PIN WWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4100 1.0200 5.8400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END WWL2

  PIN WBL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8400 1.0500 2.3850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1872 ;
  END WBL1

  PIN WBL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.1300 1.0500 6.5700 1.1500 ;
    END
    ANTENNAGATEAREA 0.1872 ;
  END WBL2

  PIN WWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.7750 4.1500 1.4900 ;
        RECT 3.4000 0.6850 4.1500 0.7750 ;
        RECT 3.4000 0.7750 3.4900 1.0100 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END WWL1

  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9600 0.3500 1.3500 ;
        RECT 0.2500 1.3500 0.4300 1.4400 ;
        RECT 0.2500 0.8700 0.4300 0.9600 ;
        RECT 0.3400 1.4400 0.4300 1.7400 ;
        RECT 0.3400 0.5900 0.4300 0.8700 ;
    END
    ANTENNADIFFAREA 0.286 ;
  END RBL1

  PIN RBL2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.4500 0.9250 8.5500 1.4350 ;
        RECT 8.4300 1.4350 8.5500 1.8050 ;
        RECT 8.4300 0.5700 8.5500 0.9250 ;
        RECT 7.9100 0.4800 8.5500 0.5700 ;
        RECT 7.9100 0.5700 8.0100 1.6850 ;
    END
    ANTENNADIFFAREA 0.4576 ;
  END RBL2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.6450 2.7200 ;
        RECT 4.8600 2.0100 5.0700 2.0800 ;
        RECT 6.2000 2.0100 6.2900 2.0800 ;
        RECT 6.8150 2.0100 6.9050 2.0800 ;
        RECT 7.3600 2.0100 7.4500 2.0800 ;
        RECT 2.2450 1.9600 2.3350 2.0800 ;
        RECT 1.7250 1.8900 1.8150 2.0800 ;
        RECT 4.3600 1.8500 4.5700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8500 1.3250 0.9400 1.7250 ;
      RECT 0.7800 1.1150 0.9400 1.3250 ;
      RECT 0.8500 0.4700 0.9400 1.1150 ;
      RECT 0.0700 1.8300 1.5400 1.9200 ;
      RECT 1.4500 0.5500 1.5400 1.8300 ;
      RECT 0.6000 0.5400 0.6900 1.8300 ;
      RECT 0.0700 1.5300 0.1700 1.8300 ;
      RECT 0.0700 0.7800 0.1600 1.5300 ;
      RECT 0.0700 0.4100 0.1700 0.7800 ;
      RECT 2.9350 1.3500 3.1650 1.4400 ;
      RECT 2.9350 1.0300 3.0250 1.3500 ;
      RECT 2.9350 0.9400 3.1050 1.0300 ;
      RECT 3.0150 0.5700 3.1050 0.9400 ;
      RECT 2.4950 0.4800 3.1050 0.5700 ;
      RECT 2.4950 0.5700 2.5850 0.7600 ;
      RECT 1.9850 0.7600 2.5850 0.8500 ;
      RECT 2.4950 0.8500 2.5850 1.2450 ;
      RECT 1.9850 1.2450 2.5850 1.3350 ;
      RECT 2.4950 1.3350 2.5850 1.6200 ;
      RECT 1.9850 0.4800 2.0750 0.7600 ;
      RECT 1.9850 1.3350 2.0750 1.6200 ;
      RECT 3.1150 1.1400 3.7800 1.2300 ;
      RECT 3.2350 1.5300 3.4450 1.6200 ;
      RECT 3.3550 1.2300 3.4450 1.5300 ;
      RECT 3.2200 0.4100 3.3100 1.1400 ;
      RECT 4.5250 1.1800 4.6150 1.5800 ;
      RECT 4.3000 1.0700 4.6150 1.1800 ;
      RECT 4.5250 0.8300 4.6150 1.0700 ;
      RECT 4.5250 0.7400 4.7750 0.8300 ;
      RECT 5.1800 1.2600 5.8400 1.3500 ;
      RECT 5.1800 1.3500 5.2700 1.7400 ;
      RECT 5.1800 0.5950 5.2700 1.2600 ;
      RECT 3.8350 0.5050 5.2700 0.5950 ;
      RECT 5.1800 0.4850 5.2700 0.5050 ;
      RECT 3.8350 0.4100 4.0250 0.5050 ;
      RECT 5.4300 1.4400 6.5500 1.5300 ;
      RECT 6.4600 1.5300 6.5500 1.7400 ;
      RECT 6.4600 1.3700 6.5500 1.4400 ;
      RECT 5.9500 0.6600 6.5500 0.7500 ;
      RECT 6.4600 0.7500 6.5500 0.8750 ;
      RECT 5.4300 1.5300 5.5200 1.7400 ;
      RECT 5.9500 1.5300 6.0400 1.7400 ;
      RECT 5.9500 0.9300 6.0400 1.4400 ;
      RECT 5.4300 0.8400 6.0400 0.9300 ;
      RECT 5.9500 0.7500 6.0400 0.8400 ;
      RECT 5.4300 0.5000 5.5200 0.8400 ;
      RECT 6.6600 1.0500 7.0100 1.2200 ;
      RECT 1.6500 1.0300 1.7400 1.7100 ;
      RECT 2.7550 0.6600 2.8450 1.7100 ;
      RECT 4.7200 1.8300 6.7500 1.9200 ;
      RECT 6.6600 1.2200 6.7500 1.8300 ;
      RECT 6.6600 0.5700 6.7500 1.0500 ;
      RECT 5.6900 0.4800 6.7500 0.5700 ;
      RECT 5.6900 1.9200 5.7800 1.9900 ;
      RECT 5.6900 1.6200 5.7800 1.8300 ;
      RECT 5.6900 0.5700 5.7800 0.7250 ;
      RECT 4.7200 1.7600 4.8200 1.8300 ;
      RECT 1.6500 1.7100 4.8200 1.7600 ;
      RECT 3.8700 1.6700 4.8200 1.7100 ;
      RECT 4.7300 1.0700 4.8200 1.6700 ;
      RECT 1.6500 1.7600 3.9600 1.8000 ;
      RECT 3.7600 1.8000 3.9600 1.8400 ;
      RECT 3.8700 0.9550 3.9600 1.6700 ;
      RECT 3.7600 1.8400 3.8500 1.9900 ;
      RECT 3.6000 0.8650 3.9600 0.9550 ;
      RECT 7.6600 1.4050 7.7500 1.6800 ;
      RECT 7.6600 1.1950 7.8200 1.4050 ;
      RECT 7.6600 0.5550 7.7500 1.1950 ;
      RECT 7.1000 1.8300 8.2600 1.9200 ;
      RECT 8.1700 0.6600 8.2600 1.8300 ;
      RECT 7.1000 0.5700 7.1900 1.8300 ;
  END
END RF2R2WS_X2M_A12TH

MACRO SDFFNQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.9500 0.3200 1.0500 0.6400 ;
        RECT 3.9950 0.3200 4.1650 0.4400 ;
        RECT 4.9050 0.3200 5.0050 0.6700 ;
    END
  END VSS

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5450 0.9900 4.7500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END CKN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0700 0.4050 1.4400 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 1.3100 4.3850 1.6800 ;
        RECT 4.2500 0.8600 4.3500 1.3100 ;
        RECT 4.2500 0.7700 4.4450 0.8600 ;
    END
    ANTENNADIFFAREA 0.273875 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0600 0.9700 1.4300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 0.9900 1.8050 1.1000 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.1600 1.4800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3150 1.8850 0.7300 1.9700 ;
      RECT 0.0600 1.8700 0.7300 1.8850 ;
      RECT 0.0600 1.7850 0.4150 1.8700 ;
      RECT 0.0600 0.5700 0.7600 0.6700 ;
      RECT 0.6600 0.5250 0.7600 0.5700 ;
      RECT 0.6600 0.4250 0.8300 0.5250 ;
      RECT 0.0600 0.6700 0.1600 1.7850 ;
      RECT 0.4750 1.5250 1.5400 1.6350 ;
      RECT 1.4500 1.6350 1.5400 1.9250 ;
      RECT 0.4250 0.8550 1.5550 0.9550 ;
      RECT 1.4450 0.7550 1.5550 0.8550 ;
      RECT 1.0600 0.9550 1.1600 1.5250 ;
      RECT 0.4750 1.6350 0.5800 1.7000 ;
      RECT 1.6700 1.5700 1.9150 1.6600 ;
      RECT 1.8250 0.7800 1.9150 1.5700 ;
      RECT 1.8250 0.6900 2.4800 0.7800 ;
      RECT 2.3900 0.7800 2.4800 1.2350 ;
      RECT 2.1400 1.5850 2.6600 1.6750 ;
      RECT 2.1400 1.1600 2.2300 1.5850 ;
      RECT 2.5700 0.8100 2.6600 1.5850 ;
      RECT 2.5700 0.7200 2.8300 0.8100 ;
      RECT 2.8300 1.6150 3.0350 1.7050 ;
      RECT 2.9450 0.8150 3.0350 1.6150 ;
      RECT 2.9450 0.7150 3.4850 0.8150 ;
      RECT 3.3850 0.8150 3.4850 1.0800 ;
      RECT 3.3850 1.0800 3.7800 1.1800 ;
      RECT 3.3250 1.6100 3.9600 1.7000 ;
      RECT 3.3250 1.3100 3.4150 1.6100 ;
      RECT 3.8700 1.1700 3.9600 1.6100 ;
      RECT 3.8700 1.0800 4.1400 1.1700 ;
      RECT 3.8700 0.9100 3.9600 1.0800 ;
      RECT 3.7700 0.8200 3.9600 0.9100 ;
      RECT 4.5750 1.3450 5.0700 1.4350 ;
      RECT 4.9800 0.8700 5.0700 1.3450 ;
      RECT 4.5750 0.7800 5.0700 0.8700 ;
      RECT 1.6450 0.4800 3.6850 0.5700 ;
      RECT 1.6450 0.5700 1.7350 1.4350 ;
      RECT 1.8550 0.4300 2.0550 0.4800 ;
      RECT 2.7800 0.4150 3.0100 0.4800 ;
      RECT 4.5750 1.4350 4.6650 1.7150 ;
      RECT 4.5750 0.6600 4.6650 0.7800 ;
      RECT 3.5950 0.5700 4.6650 0.6600 ;
      RECT 1.8150 1.8200 5.3200 1.9200 ;
      RECT 5.2200 0.7150 5.3200 1.8200 ;
      RECT 2.7150 1.9200 2.8850 1.9900 ;
      RECT 3.1350 0.9550 3.2250 1.8200 ;
  END
END SDFFNQ_X1M_A12TH

MACRO SDFFNQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.9850 0.3200 1.0850 0.7650 ;
        RECT 3.3600 0.3200 3.6500 0.3850 ;
        RECT 4.0000 0.3200 4.1700 0.4700 ;
        RECT 4.5350 0.3200 4.8700 0.4700 ;
        RECT 5.1050 0.3200 5.5150 0.3650 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0700 0.4050 1.4400 ;
    END
    ANTENNAGATEAREA 0.0837 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2450 1.3100 4.3900 1.6800 ;
        RECT 4.2450 0.8350 4.3450 1.3100 ;
        RECT 4.2450 0.7450 4.4500 0.8350 ;
    END
    ANTENNADIFFAREA 0.301 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0600 0.9700 1.4300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 4.5600 2.0400 4.8500 2.0800 ;
        RECT 2.1950 2.0350 2.3650 2.0800 ;
        RECT 3.3700 2.0300 3.6600 2.0800 ;
        RECT 0.9800 1.8400 1.0900 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.2100 1.4650 1.3900 ;
        RECT 1.3750 1.0550 1.4650 1.2100 ;
    END
    ANTENNAGATEAREA 0.0714 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6250 1.0500 5.0450 1.1500 ;
    END
    ANTENNAGATEAREA 0.0369 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.3100 1.8850 0.7200 1.9650 ;
      RECT 0.0600 1.8650 0.7200 1.8850 ;
      RECT 0.0600 1.7850 0.4100 1.8650 ;
      RECT 0.0600 0.5700 0.7100 0.6700 ;
      RECT 0.6100 0.5250 0.7100 0.5700 ;
      RECT 0.6100 0.4250 0.8200 0.5250 ;
      RECT 0.0600 0.6700 0.1600 1.7850 ;
      RECT 0.4750 1.5250 1.5400 1.6350 ;
      RECT 1.4500 1.6350 1.5400 1.9150 ;
      RECT 0.4050 0.8550 1.5600 0.9550 ;
      RECT 1.4700 0.6900 1.5600 0.8550 ;
      RECT 1.0600 0.9550 1.1600 1.5250 ;
      RECT 0.4750 1.6350 0.5800 1.7000 ;
      RECT 1.6600 1.5500 1.9200 1.6400 ;
      RECT 1.8300 0.7800 1.9200 1.5500 ;
      RECT 1.8300 0.6900 2.4850 0.7800 ;
      RECT 2.3950 0.7800 2.4850 1.2250 ;
      RECT 2.1400 1.5850 2.6650 1.6750 ;
      RECT 2.1400 1.1450 2.2300 1.5850 ;
      RECT 2.5750 0.8600 2.6650 1.5850 ;
      RECT 2.5750 0.7700 2.8500 0.8600 ;
      RECT 3.6750 1.1000 3.7750 1.4100 ;
      RECT 3.3900 1.0000 3.7750 1.1000 ;
      RECT 3.3900 0.8150 3.4900 1.0000 ;
      RECT 2.9500 0.7150 3.4900 0.8150 ;
      RECT 2.9500 0.8150 3.0400 1.6950 ;
      RECT 3.3550 1.6100 3.9650 1.7000 ;
      RECT 3.3550 1.2250 3.4450 1.6100 ;
      RECT 3.8750 1.1700 3.9650 1.6100 ;
      RECT 3.8750 1.0800 4.0950 1.1700 ;
      RECT 3.8750 0.8500 3.9650 1.0800 ;
      RECT 3.7750 0.7600 3.9650 0.8500 ;
      RECT 4.8100 1.4300 4.9000 1.7100 ;
      RECT 4.8100 1.3400 5.2900 1.4300 ;
      RECT 5.2000 0.8700 5.2900 1.3400 ;
      RECT 4.8100 0.7800 5.2900 0.8700 ;
      RECT 4.8100 0.6500 4.9000 0.7800 ;
      RECT 3.6000 0.5700 4.9000 0.6500 ;
      RECT 1.6500 0.5600 4.9000 0.5700 ;
      RECT 1.6500 0.5700 1.7400 1.4350 ;
      RECT 1.6500 0.4800 3.7550 0.5600 ;
      RECT 1.8550 0.4300 2.0550 0.4800 ;
      RECT 2.7850 0.4150 3.0150 0.4800 ;
      RECT 1.8050 1.8150 5.5250 1.9150 ;
      RECT 5.4250 0.7150 5.5250 1.8150 ;
      RECT 2.7600 1.1750 2.8500 1.8150 ;
      RECT 3.1750 0.9350 3.2650 1.8150 ;
  END
END SDFFNQ_X2M_A12TH

MACRO SDFFNQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.4600 ;
        RECT 0.9900 0.3200 1.1000 0.7250 ;
        RECT 5.3150 0.3200 5.4850 0.5350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.2100 1.4750 1.3900 ;
        RECT 1.3850 1.0200 1.4750 1.2100 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0700 0.4050 1.4400 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2650 1.2500 4.8850 1.3500 ;
        RECT 4.2650 1.3500 4.3650 1.7050 ;
        RECT 4.7850 1.3500 4.8850 1.7050 ;
        RECT 4.7850 0.7600 4.8850 1.2500 ;
        RECT 4.2050 0.6600 4.8850 0.7600 ;
    END
    ANTENNADIFFAREA 0.5508 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8300 1.0600 0.9500 1.4300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 5.2800 2.0150 5.4500 2.0800 ;
        RECT 0.9850 1.7900 1.0850 2.0800 ;
    END
  END VDD

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0450 1.0000 5.2600 1.2100 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.6600 0.4150 0.8700 0.5150 ;
      RECT 0.3100 1.8850 0.7300 1.9700 ;
      RECT 0.0600 1.8700 0.7300 1.8850 ;
      RECT 0.0600 1.7850 0.4100 1.8700 ;
      RECT 0.0600 0.5700 0.7600 0.6700 ;
      RECT 0.6600 0.5150 0.7600 0.5700 ;
      RECT 0.0600 0.6700 0.1600 1.7850 ;
      RECT 1.4550 1.6500 1.5550 1.9650 ;
      RECT 0.4300 1.5600 1.5550 1.6500 ;
      RECT 0.4100 0.8200 1.5500 0.9200 ;
      RECT 1.4500 0.6400 1.5500 0.8200 ;
      RECT 1.0400 0.9200 1.1400 1.5600 ;
      RECT 1.6650 1.5450 1.9150 1.6350 ;
      RECT 1.8250 0.7800 1.9150 1.5450 ;
      RECT 1.8250 0.6900 2.4800 0.7800 ;
      RECT 2.3900 0.7800 2.4800 1.2050 ;
      RECT 2.1400 1.5850 2.6600 1.6750 ;
      RECT 2.1400 1.1350 2.2300 1.5850 ;
      RECT 2.5700 0.8800 2.6600 1.5850 ;
      RECT 2.5700 0.7700 2.8100 0.8800 ;
      RECT 3.5300 1.0800 3.7800 1.1800 ;
      RECT 3.5300 0.8150 3.6300 1.0800 ;
      RECT 2.9450 0.7150 3.6300 0.8150 ;
      RECT 2.9450 0.8150 3.0350 1.6850 ;
      RECT 4.0150 1.0500 4.5500 1.1500 ;
      RECT 3.3400 1.6100 4.1050 1.7000 ;
      RECT 3.3400 1.2200 3.4300 1.6100 ;
      RECT 4.0150 1.1500 4.1050 1.6100 ;
      RECT 4.0150 0.9050 4.1050 1.0500 ;
      RECT 3.7450 0.8150 4.1050 0.9050 ;
      RECT 5.0350 1.4800 5.5050 1.5700 ;
      RECT 5.4150 0.7200 5.5050 1.4800 ;
      RECT 5.0400 0.6300 5.5050 0.7200 ;
      RECT 5.0350 1.5700 5.1350 1.7050 ;
      RECT 5.0400 0.5700 5.1300 0.6300 ;
      RECT 1.6450 0.4800 5.1300 0.5700 ;
      RECT 1.6450 0.5700 1.7350 1.4350 ;
      RECT 1.9000 0.4400 2.0700 0.4800 ;
      RECT 2.8000 0.4150 2.9750 0.4800 ;
      RECT 1.8050 1.8250 5.7100 1.9150 ;
      RECT 5.6100 0.4100 5.7100 1.8250 ;
      RECT 2.7500 1.2250 2.8400 1.8250 ;
      RECT 3.1600 0.9400 3.2500 1.8250 ;
  END
END SDFFNQ_X3M_A12TH

MACRO SDFFNRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4650 ;
        RECT 0.9850 0.3200 1.1550 0.7800 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0500 0.6850 1.1500 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 1.4100 5.4400 1.6500 ;
        RECT 5.3400 0.6650 5.4400 1.4100 ;
    END
    ANTENNADIFFAREA 0.2496 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.0500 3.0600 1.1500 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 2.4250 2.0650 2.5950 2.0800 ;
        RECT 4.3700 1.9400 4.5400 2.0800 ;
        RECT 1.0550 1.8000 1.1450 2.0800 ;
        RECT 5.9100 1.5000 6.0000 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9500 1.4750 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 1.0000 6.1050 1.1900 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.3500 1.8800 0.7600 1.9700 ;
      RECT 0.3500 1.8600 0.4400 1.8800 ;
      RECT 0.0550 1.7700 0.4400 1.8600 ;
      RECT 0.0550 0.6000 0.5000 0.6900 ;
      RECT 0.4100 0.5200 0.5000 0.6000 ;
      RECT 0.4100 0.4300 0.7800 0.5200 ;
      RECT 0.0550 0.6900 0.1450 1.7700 ;
      RECT 1.5200 1.7000 1.6100 1.9800 ;
      RECT 0.5050 1.6100 1.6100 1.7000 ;
      RECT 0.5050 0.8700 1.6100 0.9600 ;
      RECT 1.5200 0.7200 1.6100 0.8700 ;
      RECT 1.0600 0.9600 1.1500 1.6100 ;
      RECT 0.5050 1.4700 0.5950 1.6100 ;
      RECT 0.5050 0.7900 0.5950 0.8700 ;
      RECT 1.7200 1.6150 1.9700 1.7050 ;
      RECT 1.8800 1.1900 1.9700 1.6150 ;
      RECT 1.8800 1.1000 2.5500 1.1900 ;
      RECT 2.4500 0.9700 2.5500 1.1000 ;
      RECT 1.8800 0.7100 1.9700 1.1000 ;
      RECT 2.1850 1.5950 3.2600 1.6850 ;
      RECT 3.1700 1.1450 3.2600 1.5950 ;
      RECT 3.1700 1.0550 3.6600 1.1450 ;
      RECT 3.5700 0.9850 3.6600 1.0550 ;
      RECT 3.1700 0.8500 3.2600 1.0550 ;
      RECT 3.5700 0.8950 3.7650 0.9850 ;
      RECT 2.6650 0.7600 3.2600 0.8500 ;
      RECT 2.1850 1.3000 2.2750 1.5950 ;
      RECT 3.3600 1.5950 3.9900 1.6850 ;
      RECT 3.9000 0.8000 3.9900 1.5950 ;
      RECT 3.3700 0.7100 4.7300 0.8000 ;
      RECT 3.3700 0.8000 3.4600 0.9000 ;
      RECT 4.6400 0.8000 4.7300 1.0800 ;
      RECT 4.6400 1.0800 4.8150 1.2850 ;
      RECT 4.3750 1.5500 5.0200 1.6400 ;
      RECT 4.9300 1.1700 5.0200 1.5500 ;
      RECT 4.3750 0.9200 4.4650 1.5500 ;
      RECT 4.9300 1.0800 5.1400 1.1700 ;
      RECT 4.9300 0.7700 5.0200 1.0800 ;
      RECT 4.8400 0.6800 5.0200 0.7700 ;
      RECT 2.1050 1.8300 5.6850 1.8400 ;
      RECT 4.1300 1.7500 5.6850 1.8300 ;
      RECT 5.5950 0.7050 5.6850 1.7500 ;
      RECT 1.8750 1.8950 4.2200 1.9200 ;
      RECT 3.3550 1.9200 3.5250 1.9900 ;
      RECT 2.1050 1.8400 4.2200 1.8950 ;
      RECT 4.1300 0.9300 4.2200 1.7500 ;
      RECT 1.8750 1.9200 2.1950 1.9850 ;
      RECT 1.7000 0.4850 6.3200 0.5750 ;
      RECT 6.2300 0.5750 6.3200 1.5150 ;
      RECT 1.6550 1.3250 1.7900 1.4950 ;
      RECT 1.7000 0.5750 1.7900 1.3250 ;
  END
END SDFFNRPQ_X1M_A12TH

MACRO SDFFNRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.5450 ;
        RECT 0.9350 0.3200 1.1050 0.6850 ;
        RECT 2.8900 0.3200 3.2700 0.3900 ;
        RECT 4.1100 0.3200 4.4800 0.3850 ;
        RECT 4.9250 0.3200 5.2950 0.3800 ;
        RECT 6.2150 0.3200 6.3050 0.6100 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0450 0.6550 1.1650 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0050 2.8600 1.1450 ;
        RECT 2.6500 1.1450 2.7500 1.3850 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 2.3200 2.0450 2.4900 2.0800 ;
        RECT 0.0700 1.8900 0.1700 2.0800 ;
        RECT 0.9650 1.8400 1.0850 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.1900 1.3900 1.4400 ;
        RECT 1.2500 1.0200 1.4250 1.1900 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9550 1.2500 6.3500 1.3500 ;
        RECT 5.9550 1.3500 6.0450 1.7000 ;
        RECT 6.2500 0.8900 6.3500 1.2500 ;
        RECT 5.9500 0.7900 6.3500 0.8900 ;
        RECT 5.9500 0.4350 6.0500 0.7900 ;
    END
    ANTENNADIFFAREA 0.306 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 1.0750 0.9500 1.4450 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.0050 5.1800 1.3550 ;
    END
    ANTENNAGATEAREA 0.0369 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.2600 1.8800 0.6750 1.9700 ;
      RECT 0.2600 1.7650 0.3500 1.8800 ;
      RECT 0.0450 1.6750 0.3500 1.7650 ;
      RECT 0.0450 0.6550 0.4350 0.7450 ;
      RECT 0.3450 0.5000 0.4350 0.6550 ;
      RECT 0.3450 0.4100 0.7150 0.5000 ;
      RECT 0.0450 0.7450 0.1350 1.6750 ;
      RECT 1.4000 1.7300 1.5700 1.9700 ;
      RECT 0.4400 1.6400 1.5700 1.7300 ;
      RECT 0.4000 0.8350 1.5300 0.9250 ;
      RECT 1.4400 0.6300 1.5300 0.8350 ;
      RECT 1.0450 0.9250 1.1350 1.6400 ;
      RECT 0.4400 1.5450 0.5300 1.6400 ;
      RECT 1.6600 1.6150 1.8900 1.7050 ;
      RECT 1.8000 1.1300 1.8900 1.6150 ;
      RECT 1.8000 1.0400 2.5350 1.1300 ;
      RECT 2.4150 0.9300 2.5350 1.0400 ;
      RECT 1.8000 0.6900 1.8900 1.0400 ;
      RECT 2.1050 1.5950 3.0850 1.6850 ;
      RECT 2.9950 0.9850 3.0850 1.5950 ;
      RECT 2.9950 0.8950 3.6200 0.9850 ;
      RECT 2.9950 0.7950 3.0850 0.8950 ;
      RECT 2.5500 0.7050 3.0850 0.7950 ;
      RECT 2.1050 1.2950 2.1950 1.5950 ;
      RECT 3.1950 1.5750 3.5650 1.6650 ;
      RECT 3.4750 1.2800 3.5650 1.5750 ;
      RECT 3.4750 1.1900 3.8250 1.2800 ;
      RECT 3.7350 0.8050 3.8250 1.1900 ;
      RECT 3.2000 0.7150 4.2350 0.8050 ;
      RECT 4.1450 0.8050 4.2350 1.1250 ;
      RECT 4.1450 1.1250 4.6100 1.2150 ;
      RECT 4.3450 0.6700 5.4000 0.7600 ;
      RECT 5.3100 0.7600 5.4000 1.2100 ;
      RECT 1.6200 0.4900 4.4350 0.5800 ;
      RECT 4.3450 0.5800 4.4350 0.6700 ;
      RECT 4.8650 0.7600 4.9550 1.4700 ;
      RECT 1.5850 1.2750 1.7100 1.4450 ;
      RECT 1.6200 0.5800 1.7100 1.2750 ;
      RECT 3.6650 1.5900 5.5800 1.6800 ;
      RECT 5.4900 0.7050 5.5800 1.5900 ;
      RECT 1.8150 1.8300 3.7550 1.9200 ;
      RECT 3.3300 1.9200 3.5000 1.9700 ;
      RECT 3.6650 1.6800 3.7550 1.8300 ;
      RECT 3.9300 0.9550 4.0200 1.5900 ;
      RECT 1.8150 1.9200 1.9850 1.9700 ;
      RECT 5.7450 1.0500 6.1400 1.1500 ;
      RECT 3.8650 1.8150 5.8350 1.9050 ;
      RECT 5.7450 1.1500 5.8350 1.8150 ;
      RECT 5.7450 0.5700 5.8350 1.0500 ;
      RECT 4.5450 0.4800 5.8350 0.5700 ;
      RECT 3.8650 1.9050 3.9550 1.9850 ;
  END
END SDFFNRPQ_X2M_A12TH

MACRO SDFFNRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.5450 ;
        RECT 0.9350 0.3200 1.1050 0.6450 ;
        RECT 4.9050 0.3200 5.2750 0.3800 ;
        RECT 6.1700 0.3200 6.2600 0.6100 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0300 0.6550 1.1500 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END SE

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0050 2.8500 1.1450 ;
        RECT 2.6500 1.1450 2.7500 1.3850 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 2.3100 2.0450 2.4800 2.0800 ;
        RECT 0.0700 1.8900 0.1700 2.0800 ;
        RECT 0.9650 1.8400 1.0850 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.1900 1.3900 1.4400 ;
        RECT 1.2500 1.0200 1.4250 1.1900 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9100 1.2500 6.5250 1.3500 ;
        RECT 5.9100 1.3500 6.0000 1.7000 ;
        RECT 6.4250 1.3500 6.5250 1.7000 ;
        RECT 6.4250 0.8900 6.5250 1.2500 ;
        RECT 5.9050 0.7900 6.5250 0.8900 ;
        RECT 5.9050 0.4350 6.0050 0.7900 ;
        RECT 6.4250 0.4350 6.5250 0.7900 ;
    END
    ANTENNADIFFAREA 0.5544 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 1.0750 0.9500 1.4450 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0350 1.0050 5.1650 1.3550 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.2600 1.8800 0.6750 1.9700 ;
      RECT 0.2600 1.7650 0.3500 1.8800 ;
      RECT 0.0450 1.6750 0.3500 1.7650 ;
      RECT 0.0450 0.6350 0.4350 0.7250 ;
      RECT 0.3450 0.5000 0.4350 0.6350 ;
      RECT 0.3450 0.4100 0.7150 0.5000 ;
      RECT 0.0450 0.7250 0.1350 1.6750 ;
      RECT 1.4000 1.7300 1.5700 1.9700 ;
      RECT 0.4400 1.6400 1.5700 1.7300 ;
      RECT 0.4000 0.8150 1.5300 0.9050 ;
      RECT 1.4400 0.6550 1.5300 0.8150 ;
      RECT 1.0450 0.9050 1.1350 1.6400 ;
      RECT 0.4400 1.5450 0.5300 1.6400 ;
      RECT 1.6600 1.6150 1.8900 1.7050 ;
      RECT 1.8000 1.1300 1.8900 1.6150 ;
      RECT 1.8000 1.0400 2.5250 1.1300 ;
      RECT 2.4050 0.9300 2.5250 1.0400 ;
      RECT 1.8000 0.6900 1.8900 1.0400 ;
      RECT 2.1050 1.5950 3.0750 1.6850 ;
      RECT 2.9850 0.9900 3.0750 1.5950 ;
      RECT 2.9850 0.9000 3.6100 0.9900 ;
      RECT 2.9850 0.7950 3.0750 0.9000 ;
      RECT 2.5400 0.7050 3.0750 0.7950 ;
      RECT 2.1050 1.2950 2.1950 1.5950 ;
      RECT 3.1850 1.5750 3.5550 1.6650 ;
      RECT 3.4650 1.2800 3.5550 1.5750 ;
      RECT 3.4650 1.1900 3.8150 1.2800 ;
      RECT 3.7250 0.8050 3.8150 1.1900 ;
      RECT 3.1850 0.7150 4.2150 0.8050 ;
      RECT 4.1250 0.8050 4.2150 1.1250 ;
      RECT 4.1250 1.1250 4.5900 1.2150 ;
      RECT 4.3250 0.6700 5.3550 0.7600 ;
      RECT 5.2650 0.7600 5.3550 1.2100 ;
      RECT 1.6200 0.4900 4.4150 0.5800 ;
      RECT 4.3250 0.5800 4.4150 0.6700 ;
      RECT 4.8450 0.7600 4.9350 1.4700 ;
      RECT 1.5850 1.2750 1.7100 1.4450 ;
      RECT 1.6200 0.5800 1.7100 1.2750 ;
      RECT 3.6550 1.5900 5.5350 1.6800 ;
      RECT 5.4450 0.7050 5.5350 1.5900 ;
      RECT 1.8150 1.8300 3.7450 1.9200 ;
      RECT 3.3200 1.9200 3.4900 1.9700 ;
      RECT 3.6550 1.6800 3.7450 1.8300 ;
      RECT 3.9200 0.9400 4.0100 1.5900 ;
      RECT 1.8150 1.9200 1.9850 1.9700 ;
      RECT 5.7100 1.0500 6.2050 1.1500 ;
      RECT 3.8550 1.8150 5.8000 1.9050 ;
      RECT 5.7100 1.1500 5.8000 1.8150 ;
      RECT 5.7100 0.5700 5.8000 1.0500 ;
      RECT 4.5250 0.4800 5.8000 0.5700 ;
      RECT 3.8550 1.9050 3.9450 1.9850 ;
  END
END SDFFNRPQ_X3M_A12TH

MACRO SDFFNSQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.9200 ;
        RECT 1.0950 0.3200 1.2650 0.7900 ;
        RECT 2.5600 0.3200 2.7300 0.7050 ;
        RECT 4.2100 0.3200 4.4200 0.5350 ;
        RECT 4.8050 0.3200 5.0150 0.4650 ;
        RECT 5.7150 0.3200 5.8850 0.4800 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.9100 5.1500 1.2600 ;
        RECT 5.0500 1.2600 5.2150 1.4100 ;
        RECT 5.0500 0.8100 5.2750 0.9100 ;
        RECT 5.1250 1.4100 5.2150 1.6700 ;
    END
    ANTENNADIFFAREA 0.2448 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.8100 2.0100 3.0200 2.0800 ;
        RECT 1.0650 1.8800 1.2350 2.0800 ;
        RECT 0.0850 1.6800 0.1850 2.0800 ;
        RECT 5.7050 1.6800 5.7950 2.0800 ;
    END
  END VDD

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.1650 5.7500 1.4950 ;
        RECT 5.6500 1.0750 5.9050 1.1650 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END CKN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1700 1.5050 ;
    END
    ANTENNAGATEAREA 0.0684 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0300 1.0600 1.1500 1.4500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0800 1.5700 1.5150 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6900 1.4500 3.0450 1.5500 ;
        RECT 2.9450 1.1950 3.0450 1.4500 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END SN
  OBS
    LAYER M1 ;
      RECT 0.3450 1.8800 0.7200 1.9700 ;
      RECT 0.3450 0.5900 0.4450 1.8800 ;
      RECT 0.3450 0.4900 0.6700 0.5900 ;
      RECT 1.5450 1.7700 1.7150 1.9700 ;
      RECT 0.5950 1.6800 1.7150 1.7700 ;
      RECT 0.5950 0.8800 1.6750 0.9700 ;
      RECT 1.5850 0.7550 1.6750 0.8800 ;
      RECT 0.5950 0.9700 0.6850 1.6800 ;
      RECT 0.5950 0.7550 0.6850 0.8800 ;
      RECT 1.8050 1.5950 2.0800 1.6850 ;
      RECT 1.9900 1.1700 2.0800 1.5950 ;
      RECT 1.9900 1.0800 2.6800 1.1700 ;
      RECT 2.5900 1.1700 2.6800 1.2900 ;
      RECT 1.9900 0.7450 2.0800 1.0800 ;
      RECT 2.2500 1.6400 3.2350 1.7400 ;
      RECT 3.1350 0.7550 3.2350 1.6400 ;
      RECT 2.2500 1.2900 2.3500 1.6400 ;
      RECT 3.3750 1.6500 4.3750 1.7400 ;
      RECT 4.2850 1.1700 4.3750 1.6500 ;
      RECT 3.3750 0.9650 3.4650 1.6500 ;
      RECT 4.2850 1.0800 4.7400 1.1700 ;
      RECT 3.3750 0.7550 3.5200 0.9650 ;
      RECT 4.5350 1.4150 4.6250 1.7400 ;
      RECT 4.5350 1.3250 4.9600 1.4150 ;
      RECT 4.8700 0.9350 4.9600 1.3250 ;
      RECT 3.8200 0.8450 4.9600 0.9350 ;
      RECT 3.8200 0.9350 3.9100 1.5350 ;
      RECT 1.9150 1.8300 5.4800 1.9200 ;
      RECT 5.3900 0.7500 5.4800 1.8300 ;
      RECT 3.2600 1.9200 3.4700 1.9900 ;
      RECT 1.9150 1.9200 2.1250 1.9600 ;
      RECT 3.6100 0.6350 6.1200 0.6600 ;
      RECT 6.0300 0.6600 6.1200 1.5550 ;
      RECT 4.6150 0.5700 6.1200 0.6350 ;
      RECT 2.3500 0.6050 2.4400 0.8550 ;
      RECT 1.7800 0.5150 2.4400 0.6050 ;
      RECT 1.7800 0.6050 1.8700 1.3500 ;
      RECT 1.6800 1.3500 1.8700 1.4400 ;
      RECT 3.5800 1.3650 3.7000 1.5500 ;
      RECT 3.6100 0.7250 3.7000 1.3650 ;
      RECT 3.6100 0.5700 3.7000 0.6350 ;
      RECT 2.8500 0.4800 3.7000 0.5700 ;
      RECT 3.2950 0.4350 3.5050 0.4800 ;
      RECT 2.8500 0.5700 2.9400 0.8550 ;
      RECT 2.3500 0.8550 2.9400 0.9450 ;
      RECT 3.6100 0.6600 4.7050 0.7250 ;
      RECT 5.3850 0.5000 5.5950 0.5700 ;
  END
END SDFFNSQ_X1M_A12TH

MACRO SDFFNSQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9200 ;
        RECT 1.0500 0.3200 1.2200 0.7200 ;
        RECT 2.4900 0.3200 2.5900 0.4300 ;
        RECT 5.7700 0.3200 5.8600 0.7300 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9600 2.9500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0942 ;
  END SN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8300 5.1500 1.2750 ;
        RECT 4.9450 1.2750 5.1500 1.3750 ;
        RECT 4.9450 0.6600 5.1500 0.8300 ;
        RECT 4.9450 1.3750 5.0450 1.6900 ;
    END
    ANTENNADIFFAREA 0.306 ;
  END Q

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.0804 ;
  END SE

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6100 1.0500 5.9450 1.1500 ;
        RECT 5.8550 1.1500 5.9450 1.2550 ;
    END
    ANTENNAGATEAREA 0.0369 ;
  END CKN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.7250 2.0100 2.9350 2.0800 ;
        RECT 1.0700 1.8250 1.1600 2.0800 ;
        RECT 0.0800 1.7000 0.1700 2.0800 ;
    END
  END VDD

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2900 0.9500 1.4900 ;
        RECT 0.8500 1.1200 1.0350 1.2900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 1.0650 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8300 0.8050 1.9200 ;
      RECT 0.3400 0.5500 0.4300 1.8300 ;
      RECT 0.3400 0.4600 0.6150 0.5500 ;
      RECT 1.5300 1.7050 1.6200 1.9850 ;
      RECT 0.5700 1.6150 1.6200 1.7050 ;
      RECT 0.5700 0.8100 1.6300 0.9000 ;
      RECT 1.5400 0.6650 1.6300 0.8100 ;
      RECT 0.5700 0.9000 0.6600 1.6150 ;
      RECT 0.5700 0.6950 0.6600 0.8100 ;
      RECT 1.7300 1.5400 2.0250 1.6300 ;
      RECT 1.9350 0.8450 2.0250 1.5400 ;
      RECT 1.9350 0.7550 2.7200 0.8450 ;
      RECT 2.6300 0.8450 2.7200 1.3850 ;
      RECT 2.2150 1.6500 3.1350 1.7400 ;
      RECT 3.0450 0.8100 3.1350 1.6500 ;
      RECT 2.9200 0.7200 3.1350 0.8100 ;
      RECT 2.2150 1.1800 2.3050 1.6500 ;
      RECT 3.2550 1.5800 4.2500 1.6700 ;
      RECT 3.2550 1.5250 3.4400 1.5800 ;
      RECT 4.1600 1.1350 4.2500 1.5800 ;
      RECT 3.2550 0.6800 3.3450 1.5250 ;
      RECT 4.1600 1.0450 4.5650 1.1350 ;
      RECT 4.3900 1.4150 4.4800 1.7150 ;
      RECT 4.3900 1.3250 4.8450 1.4150 ;
      RECT 4.7550 0.8000 4.8450 1.3250 ;
      RECT 3.7250 0.7100 4.8450 0.8000 ;
      RECT 3.7250 0.8000 3.8150 1.3050 ;
      RECT 1.8600 1.8300 5.5000 1.9200 ;
      RECT 5.4100 0.6800 5.5000 1.8300 ;
      RECT 3.4300 1.9200 3.6400 1.9900 ;
      RECT 6.0300 1.4900 6.1200 1.7900 ;
      RECT 6.0300 1.4000 6.1550 1.4900 ;
      RECT 6.0650 0.9300 6.1550 1.4000 ;
      RECT 5.5900 0.8400 6.1550 0.9300 ;
      RECT 6.0300 0.5750 6.1550 0.8400 ;
      RECT 2.0100 0.5250 2.1800 0.5350 ;
      RECT 1.7250 0.6250 1.8150 1.2200 ;
      RECT 1.6750 1.2200 1.8150 1.4100 ;
      RECT 3.5350 0.5700 3.6250 1.2400 ;
      RECT 3.4550 1.2400 3.6250 1.3300 ;
      RECT 1.7250 0.5700 2.8200 0.6250 ;
      RECT 5.5900 0.5700 5.6800 0.8400 ;
      RECT 1.7250 0.5350 5.6800 0.5700 ;
      RECT 2.7300 0.4800 5.6800 0.5350 ;
      RECT 5.4450 0.4200 5.6800 0.4800 ;
  END
END SDFFNSQ_X2M_A12TH

MACRO SDFFNSQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.9200 ;
        RECT 1.0500 0.3200 1.2200 0.6300 ;
        RECT 4.2600 0.3200 4.3600 0.5100 ;
        RECT 4.7650 0.3200 4.9350 0.5000 ;
        RECT 5.2850 0.3200 5.4550 0.5000 ;
        RECT 6.1100 0.3200 6.2800 0.5350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 3.9300 2.0200 4.1400 2.0800 ;
        RECT 2.7650 2.0100 2.9750 2.0800 ;
        RECT 1.0850 1.8000 1.1850 2.0800 ;
        RECT 0.0850 1.6800 0.1850 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 0.9750 1.5550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.0500 1.2100 1.1500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.8600 5.9500 1.2800 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END CKN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0600 1.2500 5.6800 1.3500 ;
        RECT 5.0600 1.3500 5.1600 1.6900 ;
        RECT 5.5800 1.3500 5.6800 1.6900 ;
        RECT 5.5800 0.9100 5.6800 1.2500 ;
        RECT 5.0250 0.8100 5.6800 0.9100 ;
    END
    ANTENNADIFFAREA 0.5601 ;
  END Q

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0300 3.0100 1.4150 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END SN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.3450 1.7750 0.7850 1.8750 ;
      RECT 0.3450 0.5300 0.4450 1.7750 ;
      RECT 0.3450 0.4300 0.6250 0.5300 ;
      RECT 1.5450 1.6000 1.6450 1.9200 ;
      RECT 0.5400 1.5100 1.6450 1.6000 ;
      RECT 0.5400 0.7500 1.6500 0.8400 ;
      RECT 1.5600 0.6400 1.6500 0.7500 ;
      RECT 0.5400 0.8400 0.6300 1.5100 ;
      RECT 1.7600 1.5150 2.0400 1.6050 ;
      RECT 1.9500 0.8400 2.0400 1.5150 ;
      RECT 1.9500 0.7500 2.7200 0.8400 ;
      RECT 2.6300 0.8400 2.7200 1.3150 ;
      RECT 2.2500 1.6100 3.2350 1.7100 ;
      RECT 3.1350 0.8050 3.2350 1.6100 ;
      RECT 2.9900 0.7050 3.2350 0.8050 ;
      RECT 2.2500 1.1800 2.3500 1.6100 ;
      RECT 3.3500 1.4650 4.4350 1.5550 ;
      RECT 4.3450 1.1600 4.4350 1.4650 ;
      RECT 3.3500 0.7250 3.4400 1.4650 ;
      RECT 4.3450 1.0600 4.7400 1.1600 ;
      RECT 4.8350 1.0500 5.3400 1.1500 ;
      RECT 4.5400 1.3750 4.6400 1.6500 ;
      RECT 4.5400 1.2750 4.9250 1.3750 ;
      RECT 4.8350 1.1500 4.9250 1.2750 ;
      RECT 4.8350 0.9250 4.9250 1.0500 ;
      RECT 3.8600 0.8250 4.9250 0.9250 ;
      RECT 3.8600 0.9250 3.9600 1.3650 ;
      RECT 5.8050 1.4200 6.3250 1.5100 ;
      RECT 6.2350 0.7350 6.3250 1.4200 ;
      RECT 5.8550 0.7000 6.3250 0.7350 ;
      RECT 3.5850 0.6450 6.3250 0.7000 ;
      RECT 3.5850 0.7000 3.6750 1.3700 ;
      RECT 3.5850 0.5700 3.6750 0.6100 ;
      RECT 1.7400 0.4800 3.6750 0.5700 ;
      RECT 3.3750 0.4100 3.5450 0.4800 ;
      RECT 1.7400 0.5700 1.8300 1.4050 ;
      RECT 3.5850 0.6100 5.9650 0.6450 ;
      RECT 5.8550 0.5000 5.9650 0.6100 ;
      RECT 5.8850 1.6550 6.5050 1.7450 ;
      RECT 6.4150 0.4100 6.5050 1.6550 ;
      RECT 3.4900 1.9200 3.7000 1.9750 ;
      RECT 1.8850 1.9200 2.0950 1.9550 ;
      RECT 1.8850 1.8300 5.9750 1.9200 ;
      RECT 5.8850 1.7450 5.9750 1.8300 ;
  END
END SDFFNSQ_X3M_A12TH

MACRO SDFFNSRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.0750 0.3200 0.2150 0.4650 ;
        RECT 0.9700 0.3200 1.0700 0.7200 ;
        RECT 3.7750 0.3200 4.1850 0.3700 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.4100 1.5050 ;
    END
    ANTENNAGATEAREA 0.0648 ;
  END SE

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0950 4.2500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0873 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 1.1900 5.3500 1.5000 ;
        RECT 5.0950 1.0900 5.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0753 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 1.2900 6.2450 1.6800 ;
        RECT 6.0500 0.8300 6.1500 1.2900 ;
        RECT 6.0500 0.6600 6.2450 0.8300 ;
    END
    ANTENNADIFFAREA 0.2464 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 2.3450 1.9650 2.5150 2.0800 ;
        RECT 3.2100 1.9650 3.3800 2.0800 ;
        RECT 1.0000 1.8300 1.1700 2.0800 ;
        RECT 6.7500 1.7000 6.8500 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0800 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0550 0.9600 1.5000 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 1.2100 6.9250 1.3800 ;
        RECT 6.6500 1.3800 6.7500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 6.5500 1.0000 7.1050 1.0900 ;
      RECT 7.0150 1.0900 7.1050 1.7350 ;
      RECT 7.0150 0.7050 7.1050 1.0000 ;
      RECT 1.6800 0.4800 6.6400 0.5700 ;
      RECT 6.5500 0.5700 6.6400 1.0000 ;
      RECT 4.4000 0.5700 4.4900 1.5350 ;
      RECT 1.6600 1.3000 1.7700 1.4700 ;
      RECT 1.6800 0.5700 1.7700 1.3000 ;
      RECT 0.3800 1.9000 0.7500 1.9900 ;
      RECT 0.3800 1.8750 0.4700 1.9000 ;
      RECT 0.0600 1.7850 0.4700 1.8750 ;
      RECT 0.0600 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5100 0.5100 0.6000 ;
      RECT 0.4200 0.4200 0.7950 0.5100 ;
      RECT 0.0600 0.6900 0.1500 1.7850 ;
      RECT 1.4600 1.7200 1.6300 1.9500 ;
      RECT 0.6700 1.6850 1.6300 1.7200 ;
      RECT 0.4550 1.6300 1.6300 1.6850 ;
      RECT 0.3850 0.8300 1.5900 0.9200 ;
      RECT 1.5000 0.6700 1.5900 0.8300 ;
      RECT 1.1450 0.9200 1.2350 1.6300 ;
      RECT 0.4550 1.5950 0.7600 1.6300 ;
      RECT 1.7250 1.5900 1.9500 1.6800 ;
      RECT 1.8600 1.1900 1.9500 1.5900 ;
      RECT 1.8600 1.1000 2.9200 1.1900 ;
      RECT 2.8300 1.1900 2.9200 1.4600 ;
      RECT 1.8600 0.6800 1.9500 1.1000 ;
      RECT 2.6700 0.6700 3.3900 0.7600 ;
      RECT 2.1700 1.5700 3.5900 1.6600 ;
      RECT 2.1700 1.3050 2.2600 1.5700 ;
      RECT 3.4800 0.9550 3.5900 1.5700 ;
      RECT 2.9300 0.8650 3.5900 0.9550 ;
      RECT 3.5000 0.7050 3.5900 0.8650 ;
      RECT 4.5900 0.6700 5.5850 0.7600 ;
      RECT 5.4950 0.7600 5.5850 1.2700 ;
      RECT 3.7400 1.6450 4.6800 1.7350 ;
      RECT 4.5900 0.7600 4.6800 1.6450 ;
      RECT 3.7400 0.6950 3.8500 1.6450 ;
      RECT 4.9800 1.6400 5.8500 1.7300 ;
      RECT 5.7600 1.1950 5.8500 1.6400 ;
      RECT 5.7600 1.0250 5.9250 1.1950 ;
      RECT 5.7600 0.8850 5.8500 1.0250 ;
      RECT 5.6750 0.6950 5.8500 0.8850 ;
      RECT 4.9800 1.3500 5.0700 1.6400 ;
      RECT 3.4950 1.8600 6.5200 1.9200 ;
      RECT 1.8600 1.8300 6.5200 1.8600 ;
      RECT 6.3700 1.5550 6.5200 1.8300 ;
      RECT 6.3700 0.6850 6.4600 1.5550 ;
      RECT 4.7900 0.8850 4.8800 1.8300 ;
      RECT 3.4950 1.9200 3.8150 1.9700 ;
      RECT 2.0350 1.7700 3.5900 1.8300 ;
      RECT 1.8600 1.8600 2.1250 1.9200 ;
  END
END SDFFNSRPQ_X1M_A12TH

MACRO SDFFNSRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.4850 ;
        RECT 0.9900 0.3200 1.0900 0.7250 ;
        RECT 6.9650 0.3200 7.0650 0.7300 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.3700 1.5000 ;
    END
    ANTENNAGATEAREA 0.0792 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8200 1.0350 0.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1450 4.1700 1.5100 ;
    END
    ANTENNAGATEAREA 0.1014 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1450 1.0100 5.3500 1.4550 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 1.2900 6.2050 1.7150 ;
        RECT 6.0500 0.7900 6.1500 1.2900 ;
        RECT 6.0500 0.6900 6.2700 0.7900 ;
    END
    ANTENNADIFFAREA 0.306 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0750 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0250 1.0700 7.1500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0369 ;
  END CKN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.4450 2.7200 ;
        RECT 5.8400 2.0400 5.9800 2.0800 ;
        RECT 2.3750 2.0250 2.5450 2.0800 ;
        RECT 5.3250 1.9850 5.4950 2.0800 ;
        RECT 0.0600 1.9450 0.2300 2.0800 ;
        RECT 3.1650 1.9200 3.2650 2.0800 ;
        RECT 6.8650 1.5100 6.9650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 7.2050 1.5150 7.3500 1.7050 ;
      RECT 7.2600 0.9300 7.3500 1.5150 ;
      RECT 6.7800 0.8400 7.3500 0.9300 ;
      RECT 7.2300 0.5900 7.3500 0.8400 ;
      RECT 6.7800 0.9300 6.8700 1.1650 ;
      RECT 6.7800 0.5700 6.8700 0.8400 ;
      RECT 1.6800 0.4800 6.8700 0.5700 ;
      RECT 4.3300 0.5700 4.4200 1.5350 ;
      RECT 1.6800 0.5700 1.7700 1.4550 ;
      RECT 0.3300 1.8800 0.7500 1.9700 ;
      RECT 0.3300 1.8350 0.4200 1.8800 ;
      RECT 0.0550 1.7450 0.4200 1.8350 ;
      RECT 0.0550 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5000 0.5100 0.6000 ;
      RECT 0.4200 0.4100 0.7950 0.5000 ;
      RECT 0.0550 0.6900 0.1450 1.7450 ;
      RECT 1.5000 1.6500 1.5900 1.9750 ;
      RECT 0.4750 1.5600 1.5900 1.6500 ;
      RECT 0.4100 0.8200 1.5900 0.9100 ;
      RECT 1.5000 0.7050 1.5900 0.8200 ;
      RECT 1.0550 0.9100 1.1450 1.5600 ;
      RECT 1.7000 1.5900 1.9500 1.6800 ;
      RECT 1.8600 1.1750 1.9500 1.5900 ;
      RECT 1.8600 1.0850 2.9200 1.1750 ;
      RECT 2.8300 1.1750 2.9200 1.2950 ;
      RECT 1.8600 0.6800 1.9500 1.0850 ;
      RECT 2.6700 0.6700 3.4000 0.7600 ;
      RECT 2.1850 1.4500 3.1350 1.5400 ;
      RECT 2.1850 1.2850 2.2750 1.4500 ;
      RECT 3.0450 0.9550 3.1350 1.4500 ;
      RECT 2.9300 0.8650 3.6050 0.9550 ;
      RECT 3.5150 0.9550 3.6050 1.3500 ;
      RECT 3.5150 0.7250 3.6050 0.8650 ;
      RECT 3.4350 1.3500 3.6050 1.5200 ;
      RECT 4.5300 0.6600 5.5600 0.7500 ;
      RECT 5.4700 0.7500 5.5600 1.3250 ;
      RECT 3.6950 1.6450 4.6200 1.7350 ;
      RECT 4.5300 0.7500 4.6200 1.6450 ;
      RECT 3.6950 1.2950 3.7850 1.6450 ;
      RECT 3.6950 1.2050 3.8800 1.2950 ;
      RECT 3.7900 0.6800 3.8800 1.2050 ;
      RECT 4.9100 1.5550 5.9450 1.6450 ;
      RECT 5.8550 1.0650 5.9450 1.5550 ;
      RECT 5.6500 0.9750 5.9450 1.0650 ;
      RECT 5.6500 0.7350 5.7400 0.9750 ;
      RECT 4.9100 1.3500 5.0000 1.5550 ;
      RECT 3.4350 1.8300 6.6700 1.8600 ;
      RECT 5.5700 1.8600 6.6700 1.9200 ;
      RECT 6.5800 0.6650 6.6700 1.8300 ;
      RECT 3.4350 1.8600 5.2550 1.9200 ;
      RECT 5.1650 1.7700 5.6600 1.8300 ;
      RECT 4.7300 0.8650 4.8200 1.8300 ;
      RECT 3.4350 1.7700 3.5250 1.8300 ;
      RECT 2.1250 1.6800 3.5250 1.7700 ;
      RECT 2.1250 1.7700 2.2150 1.8300 ;
      RECT 3.2550 1.2400 3.3450 1.6800 ;
      RECT 1.9100 1.8300 2.2150 1.9200 ;
      RECT 3.2550 1.0700 3.4250 1.2400 ;
  END
END SDFFNSRPQ_X2M_A12TH

MACRO SDFFNSRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.4850 ;
        RECT 0.9900 0.3200 1.0900 0.7250 ;
        RECT 7.2800 0.3200 7.3800 0.8000 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0900 0.3700 1.5000 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8200 1.0350 0.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1450 4.1700 1.5450 ;
    END
    ANTENNAGATEAREA 0.1014 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1450 1.0100 5.3500 1.4550 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.7900 6.5500 1.2500 ;
        RECT 6.1100 1.2500 6.7300 1.3500 ;
        RECT 6.0500 0.6900 6.7850 0.7900 ;
        RECT 6.1100 1.3500 6.2100 1.7200 ;
        RECT 6.6300 1.3500 6.7300 1.7200 ;
    END
    ANTENNADIFFAREA 0.5539 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 5.8400 2.0400 5.9800 2.0800 ;
        RECT 2.3750 2.0250 2.5450 2.0800 ;
        RECT 3.1650 1.9150 3.2650 2.0800 ;
        RECT 7.1800 1.5450 7.2800 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.0200 1.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1000 1.2500 7.4550 1.3500 ;
        RECT 7.3500 1.0700 7.4550 1.2500 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 3.4350 1.8300 6.9850 1.9200 ;
      RECT 6.8950 0.7550 6.9850 1.8300 ;
      RECT 4.7300 0.8650 4.8200 1.8300 ;
      RECT 2.1250 1.6800 3.5250 1.7700 ;
      RECT 3.4350 1.7700 3.5250 1.8300 ;
      RECT 3.2550 1.2400 3.3450 1.6800 ;
      RECT 3.2550 1.0700 3.4250 1.2400 ;
      RECT 1.8650 1.8300 2.2150 1.9200 ;
      RECT 2.1250 1.7700 2.2150 1.8300 ;
      RECT 7.5400 1.6400 7.6450 1.9150 ;
      RECT 7.5400 1.5000 7.7450 1.6400 ;
      RECT 7.6550 0.9800 7.7450 1.5000 ;
      RECT 7.0800 0.8900 7.7450 0.9800 ;
      RECT 7.5450 0.6400 7.6650 0.8900 ;
      RECT 7.0800 0.5700 7.1700 0.8900 ;
      RECT 1.6800 0.4800 7.1700 0.5700 ;
      RECT 6.9000 0.4300 7.1700 0.4800 ;
      RECT 4.0150 0.5700 4.1050 1.0500 ;
      RECT 4.3300 0.5700 4.4200 1.5350 ;
      RECT 1.6800 0.5700 1.7700 1.4550 ;
      RECT 0.3300 1.8800 0.7500 1.9700 ;
      RECT 0.3300 1.7850 0.4200 1.8800 ;
      RECT 0.0550 1.6950 0.4200 1.7850 ;
      RECT 0.0550 0.6000 0.5100 0.6900 ;
      RECT 0.4200 0.5000 0.5100 0.6000 ;
      RECT 0.4200 0.4100 0.7950 0.5000 ;
      RECT 0.0550 0.6900 0.1450 1.6950 ;
      RECT 1.5000 1.7700 1.5900 1.9900 ;
      RECT 0.5150 1.6800 1.5900 1.7700 ;
      RECT 1.5000 1.6000 1.5900 1.6800 ;
      RECT 0.4100 0.8200 1.5900 0.9100 ;
      RECT 1.5000 0.7050 1.5900 0.8200 ;
      RECT 1.0550 0.9100 1.1450 1.6800 ;
      RECT 0.5150 1.5350 0.6050 1.6800 ;
      RECT 1.7250 1.5900 1.9500 1.6800 ;
      RECT 1.8600 1.1750 1.9500 1.5900 ;
      RECT 1.8600 1.0850 2.9200 1.1750 ;
      RECT 2.8300 1.1750 2.9200 1.2800 ;
      RECT 1.8600 0.6800 1.9500 1.0850 ;
      RECT 2.6700 0.6700 3.4000 0.7600 ;
      RECT 2.2100 1.4500 3.1350 1.5400 ;
      RECT 2.2100 1.2850 2.3000 1.4500 ;
      RECT 3.0450 0.9550 3.1350 1.4500 ;
      RECT 2.9300 0.8650 3.6050 0.9550 ;
      RECT 3.5150 0.9550 3.6050 1.3500 ;
      RECT 3.5150 0.6950 3.6050 0.8650 ;
      RECT 3.4350 1.3500 3.6050 1.5200 ;
      RECT 4.5300 0.6600 5.5600 0.7500 ;
      RECT 5.4700 0.7500 5.5600 1.3250 ;
      RECT 3.6950 1.6450 4.6200 1.7350 ;
      RECT 4.5300 0.7500 4.6200 1.6450 ;
      RECT 3.6950 1.2950 3.7850 1.6450 ;
      RECT 3.6950 1.2050 3.8800 1.2950 ;
      RECT 3.7900 0.7100 3.8800 1.2050 ;
      RECT 5.6500 0.9750 6.3500 1.0650 ;
      RECT 4.9100 1.5550 5.9450 1.6450 ;
      RECT 5.8550 1.0650 5.9450 1.5550 ;
      RECT 5.6500 0.7400 5.7400 0.9750 ;
      RECT 4.9100 1.3500 5.0000 1.5550 ;
  END
END SDFFNSRPQ_X3M_A12TH

MACRO SDFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7400 ;
        RECT 0.9400 0.3200 1.1100 0.4800 ;
        RECT 2.3000 0.3200 2.4000 0.7950 ;
        RECT 3.4150 0.3200 3.5150 0.6750 ;
        RECT 4.7100 0.3200 4.8100 0.5750 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.2500 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0297 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 1.0450 1.8800 1.2150 2.0800 ;
        RECT 0.3300 1.8400 0.4400 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5400 1.2100 4.7500 1.4650 ;
        RECT 4.5400 1.0750 4.6400 1.2100 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.7800 4.1600 1.2850 ;
        RECT 3.9750 1.2850 4.1600 1.4800 ;
        RECT 3.9900 0.6800 4.1600 0.7800 ;
    END
    ANTENNADIFFAREA 0.156425 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.3100 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.4500 0.8750 1.5500 ;
        RECT 0.7750 1.0050 0.8750 1.4500 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.8400 1.7650 1.7150 1.7700 ;
      RECT 1.4150 1.7700 1.7150 1.8550 ;
      RECT 0.8400 1.6800 1.5050 1.7650 ;
      RECT 0.9650 1.0100 1.5700 1.1000 ;
      RECT 1.4800 0.4300 1.5700 1.0100 ;
      RECT 0.9650 1.1000 1.0550 1.6800 ;
      RECT 0.9650 0.8500 1.0550 1.0100 ;
      RECT 0.8550 0.7500 1.0550 0.8500 ;
      RECT 0.8400 1.7700 0.9300 1.9900 ;
      RECT 1.8400 1.2650 2.6100 1.3650 ;
      RECT 2.5100 1.3650 2.6100 1.4850 ;
      RECT 1.8400 1.3650 1.9300 1.9350 ;
      RECT 1.8400 0.6800 1.9300 1.2650 ;
      RECT 2.6300 1.5950 2.8200 1.6950 ;
      RECT 2.7300 1.1750 2.8200 1.5950 ;
      RECT 2.1250 1.0850 2.8200 1.1750 ;
      RECT 2.7300 0.8500 2.8200 1.0850 ;
      RECT 2.6700 0.6800 2.8200 0.8500 ;
      RECT 2.9200 1.6100 3.6200 1.7000 ;
      RECT 3.5200 1.1850 3.6200 1.6100 ;
      RECT 2.9200 0.6800 3.0200 1.6100 ;
      RECT 3.2950 1.0750 3.3850 1.1800 ;
      RECT 3.2950 0.9850 3.8850 1.0750 ;
      RECT 3.7750 1.0750 3.8850 1.7300 ;
      RECT 3.7850 0.6800 3.8850 0.9850 ;
      RECT 2.0200 1.8300 4.9400 1.9200 ;
      RECT 4.8500 0.9750 4.9400 1.8300 ;
      RECT 4.3500 0.8850 4.9400 0.9750 ;
      RECT 4.3500 0.6800 4.4400 0.8850 ;
      RECT 2.0200 1.4750 2.1100 1.8300 ;
      RECT 4.5300 0.6850 5.1200 0.7750 ;
      RECT 5.0300 0.7750 5.1200 1.9500 ;
      RECT 2.0500 0.5700 2.1400 0.9050 ;
      RECT 1.6600 0.4800 2.1400 0.5700 ;
      RECT 1.6600 0.5700 1.7500 1.6050 ;
      RECT 2.0500 0.9050 2.5800 0.9950 ;
      RECT 2.4900 0.5700 2.5800 0.9050 ;
      RECT 2.4900 0.4800 3.2050 0.5700 ;
      RECT 3.1150 0.5700 3.2050 0.7850 ;
      RECT 3.1150 0.8750 3.2050 1.4900 ;
      RECT 3.6050 0.4800 4.6200 0.5700 ;
      RECT 4.5300 0.5700 4.6200 0.6850 ;
      RECT 3.1150 0.7850 3.6950 0.8750 ;
      RECT 3.6050 0.5700 3.6950 0.7850 ;
      RECT 0.6350 0.5700 1.2350 0.6600 ;
      RECT 1.1450 0.6600 1.2350 0.9000 ;
      RECT 0.0700 1.8150 0.2100 1.9850 ;
      RECT 0.0700 0.9200 0.1600 1.8150 ;
      RECT 0.0700 0.6850 0.1800 0.8300 ;
      RECT 0.0700 0.8300 0.7250 0.9200 ;
      RECT 0.6350 0.6600 0.7250 0.8300 ;
  END
END SDFFQN_X0P5M_A12TH

MACRO SDFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.3750 0.3200 0.4850 0.6450 ;
        RECT 2.2800 0.3200 2.3800 0.8500 ;
        RECT 4.7350 0.3200 4.8350 0.6500 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.2450 ;
        RECT 0.4500 1.2450 0.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0150 0.6650 4.1500 1.7050 ;
    END
    ANTENNADIFFAREA 0.244 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.0100 5.0250 1.1900 ;
        RECT 4.9300 1.1900 5.0250 1.4550 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 3.1550 2.0450 3.5250 2.0800 ;
        RECT 2.3150 1.9050 2.4850 2.0800 ;
        RECT 1.0700 1.8200 1.1800 2.0800 ;
        RECT 0.3350 1.6900 0.4450 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1750 1.2500 1.5350 1.3700 ;
    END
    ANTENNAGATEAREA 0.0606 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.8750 1.5500 ;
        RECT 0.7800 1.0500 0.8750 1.4500 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5550 1.2350 0.6450 ;
      RECT 1.1450 0.6450 1.2350 0.9400 ;
      RECT 0.0700 0.8050 0.7250 0.8950 ;
      RECT 0.6350 0.6450 0.7250 0.8050 ;
      RECT 0.0700 1.6950 0.2100 1.8800 ;
      RECT 0.0700 1.0000 0.1600 1.6950 ;
      RECT 0.0700 0.8950 0.2150 1.0000 ;
      RECT 1.2700 1.8750 1.6700 1.9650 ;
      RECT 1.2700 1.7300 1.3600 1.8750 ;
      RECT 0.8300 1.6400 1.3600 1.7300 ;
      RECT 0.9650 1.0500 1.5700 1.1400 ;
      RECT 1.4800 0.4300 1.5700 1.0500 ;
      RECT 0.8300 1.7300 0.9300 1.8800 ;
      RECT 0.9650 1.1400 1.0550 1.6400 ;
      RECT 0.9650 0.9250 1.0550 1.0500 ;
      RECT 0.8650 0.8100 1.0550 0.9250 ;
      RECT 1.8400 1.1600 2.5600 1.2500 ;
      RECT 1.7600 1.8700 1.9300 1.9700 ;
      RECT 1.8400 1.2500 1.9300 1.8700 ;
      RECT 1.8400 0.6800 1.9300 1.1600 ;
      RECT 2.2000 1.5450 2.7450 1.6350 ;
      RECT 2.2000 1.3450 2.2900 1.5450 ;
      RECT 2.6500 0.7650 2.7450 1.5450 ;
      RECT 2.8350 1.6500 3.6800 1.7400 ;
      RECT 3.5900 0.8850 3.6800 1.6500 ;
      RECT 2.8350 0.7800 2.9250 1.6500 ;
      RECT 2.8350 0.6800 3.0400 0.7800 ;
      RECT 3.7700 1.5500 3.9000 1.7200 ;
      RECT 3.8000 0.7750 3.9000 1.5500 ;
      RECT 3.3100 0.6750 3.9000 0.7750 ;
      RECT 3.3100 0.7750 3.4000 1.5350 ;
      RECT 2.4700 0.4800 4.5700 0.5700 ;
      RECT 4.4800 0.5700 4.5700 1.7200 ;
      RECT 3.0250 1.3850 3.2200 1.5550 ;
      RECT 3.1300 0.5700 3.2200 1.3850 ;
      RECT 2.4700 0.5700 2.5600 0.9600 ;
      RECT 2.7150 0.4100 2.8850 0.4800 ;
      RECT 2.0400 0.9600 2.5600 1.0500 ;
      RECT 2.0400 0.5700 2.1300 0.9600 ;
      RECT 1.6600 0.4800 2.1300 0.5700 ;
      RECT 1.6600 0.5700 1.7500 1.5750 ;
      RECT 4.6600 1.6650 5.1550 1.7650 ;
      RECT 4.6600 0.7600 5.1200 0.8500 ;
      RECT 5.0200 0.4500 5.1200 0.7600 ;
      RECT 2.5950 1.8300 4.7500 1.9200 ;
      RECT 4.6600 1.7650 4.7500 1.8300 ;
      RECT 4.6600 0.8500 4.7500 1.6650 ;
      RECT 2.0200 1.6100 2.1100 1.7250 ;
      RECT 2.7700 1.9200 2.9400 1.9900 ;
      RECT 2.5950 1.8150 2.6850 1.8300 ;
      RECT 2.0200 1.7250 2.6850 1.8150 ;
  END
END SDFFQN_X1M_A12TH

MACRO SDFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3300 0.3200 0.4400 0.6950 ;
        RECT 0.9950 0.3200 1.0850 0.4300 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 0.9800 5.3500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7800 4.5500 1.2900 ;
        RECT 4.3450 1.2900 4.5500 1.3900 ;
        RECT 4.2900 0.6800 4.5500 0.7800 ;
        RECT 4.3450 1.3900 4.4450 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9950 0.5900 1.4350 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 2.3750 2.0300 2.5900 2.0800 ;
        RECT 0.9400 2.0200 1.1100 2.0800 ;
        RECT 0.3300 1.7350 0.4400 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1350 1.2300 1.5450 1.3500 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.1850 0.3500 1.6050 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.0450 0.7950 0.8050 0.8850 ;
      RECT 0.7150 0.8850 0.8050 1.4850 ;
      RECT 0.0450 1.7000 0.2000 1.8950 ;
      RECT 0.0450 0.8850 0.1350 1.7000 ;
      RECT 0.0450 0.5050 0.1800 0.7950 ;
      RECT 0.7600 1.7700 1.6400 1.8700 ;
      RECT 0.7600 0.5400 1.5750 0.6300 ;
      RECT 1.4850 0.6300 1.5750 0.9550 ;
      RECT 0.9350 0.6400 1.0250 1.7700 ;
      RECT 0.7600 0.6300 1.0250 0.6400 ;
      RECT 1.7300 1.8700 1.9350 1.9700 ;
      RECT 1.8450 1.2600 1.9350 1.8700 ;
      RECT 1.8450 1.1600 2.5300 1.2600 ;
      RECT 1.8450 0.8400 1.9350 1.1600 ;
      RECT 2.7450 1.5250 2.8450 1.7400 ;
      RECT 2.1500 1.4250 2.8450 1.5250 ;
      RECT 2.6200 1.3700 2.8450 1.4250 ;
      RECT 2.6200 0.6600 2.7200 1.3700 ;
      RECT 2.9600 1.6100 3.7000 1.7000 ;
      RECT 3.6100 1.1650 3.7000 1.6100 ;
      RECT 2.9600 0.6800 3.0500 1.6100 ;
      RECT 3.6100 1.0550 3.9800 1.1650 ;
      RECT 3.8300 1.6050 4.1600 1.7050 ;
      RECT 4.0700 0.8300 4.1600 1.6050 ;
      RECT 3.3800 0.7300 4.1600 0.8300 ;
      RECT 3.3800 0.8300 3.4800 1.1800 ;
      RECT 4.8150 1.5850 5.0300 1.6850 ;
      RECT 4.8150 0.5700 4.9050 1.5850 ;
      RECT 1.6650 0.4800 4.9050 0.5700 ;
      RECT 1.6650 0.5700 1.7550 1.4950 ;
      RECT 3.1950 0.5700 3.2850 1.5100 ;
      RECT 2.7700 0.4100 2.9400 0.4800 ;
      RECT 1.5750 1.4950 1.7550 1.5950 ;
      RECT 2.0350 1.8300 5.3700 1.9200 ;
      RECT 5.2800 1.6800 5.3700 1.8300 ;
      RECT 5.2800 1.5900 5.5550 1.6800 ;
      RECT 5.4650 0.6450 5.5550 1.5900 ;
      RECT 4.9950 0.5550 5.5550 0.6450 ;
      RECT 4.9950 0.6450 5.0850 1.2900 ;
      RECT 2.8400 1.9200 3.0100 1.9900 ;
      RECT 2.0350 1.6700 2.1250 1.8300 ;
  END
END SDFFQN_X2M_A12TH

MACRO SDFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4250 ;
        RECT 0.9100 0.3200 1.0100 0.6050 ;
        RECT 4.4200 0.3200 4.6350 0.3600 ;
        RECT 5.2900 0.3200 5.4000 0.7100 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2050 0.9500 1.3900 ;
        RECT 0.7700 1.0250 0.9500 1.2050 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2200 1.2500 4.8400 1.3500 ;
        RECT 4.2200 1.3500 4.3200 1.7300 ;
        RECT 4.7400 1.3500 4.8400 1.7300 ;
        RECT 4.7400 0.7650 4.8400 1.2500 ;
        RECT 4.1850 0.6650 4.8400 0.7650 ;
    END
    ANTENNADIFFAREA 0.5544 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4450 1.0150 5.5550 1.4250 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0600 1.3950 1.3900 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0150 0.3600 1.4500 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4000 0.4200 0.7800 0.5200 ;
      RECT 0.0450 1.8200 0.7650 1.9200 ;
      RECT 0.0450 0.5700 0.5000 0.6700 ;
      RECT 0.4000 0.5200 0.5000 0.5700 ;
      RECT 0.0450 0.6700 0.1450 1.8200 ;
      RECT 1.3350 1.7300 1.5100 1.9600 ;
      RECT 0.4500 1.6400 1.5100 1.7300 ;
      RECT 0.3700 0.8100 1.4700 0.9100 ;
      RECT 1.3700 0.4650 1.4700 0.8100 ;
      RECT 0.4500 0.9100 0.5400 1.6400 ;
      RECT 1.6300 1.6400 1.9100 1.7300 ;
      RECT 1.8200 0.9800 1.9100 1.6400 ;
      RECT 1.7400 0.8750 1.9100 0.9800 ;
      RECT 1.7400 0.7850 2.4500 0.8750 ;
      RECT 2.3600 0.8750 2.4500 1.2400 ;
      RECT 2.0600 1.6150 2.6300 1.7050 ;
      RECT 2.0600 1.1600 2.1500 1.6150 ;
      RECT 2.5400 0.6850 2.6300 1.6150 ;
      RECT 3.5100 1.0900 3.9300 1.1900 ;
      RECT 3.5100 0.9100 3.6100 1.0900 ;
      RECT 2.7550 0.8100 3.6100 0.9100 ;
      RECT 2.7550 0.9100 2.8550 1.6400 ;
      RECT 3.2400 1.4700 4.1200 1.5700 ;
      RECT 3.2400 1.0300 3.3400 1.4700 ;
      RECT 4.0200 0.9450 4.1200 1.4700 ;
      RECT 3.7050 0.8450 4.1200 0.9450 ;
      RECT 1.5600 0.4800 5.0850 0.5700 ;
      RECT 4.9950 0.5700 5.0850 1.7300 ;
      RECT 1.5600 1.4100 1.7300 1.5200 ;
      RECT 1.5600 0.5700 1.6500 1.4100 ;
      RECT 2.9500 0.4100 3.1200 0.4800 ;
      RECT 1.8000 1.8200 5.7550 1.9100 ;
      RECT 5.6250 1.5350 5.7550 1.8200 ;
      RECT 5.6650 0.9000 5.7550 1.5350 ;
      RECT 5.1900 0.8100 5.7550 0.9000 ;
      RECT 5.6250 0.5100 5.7550 0.8100 ;
      RECT 5.1900 0.9000 5.2800 1.2400 ;
      RECT 1.8000 1.9100 1.9200 1.9900 ;
      RECT 2.9650 1.9100 3.2200 1.9900 ;
      RECT 2.9650 1.0000 3.0550 1.8200 ;
  END
END SDFFQN_X3M_A12TH

MACRO SDFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7400 ;
        RECT 0.9400 0.3200 1.1100 0.4800 ;
        RECT 2.3000 0.3200 2.4000 0.7950 ;
        RECT 3.4150 0.3200 3.5150 0.6750 ;
        RECT 4.7100 0.3200 4.8100 0.5750 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.2500 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 1.0450 1.8800 1.2150 2.0800 ;
        RECT 0.3300 1.8400 0.4400 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 1.2100 4.6400 1.4800 ;
        RECT 4.5400 1.0750 4.6400 1.2100 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.7800 4.1500 1.2650 ;
        RECT 3.9550 1.2650 4.1500 1.3650 ;
        RECT 3.9800 0.6800 4.1500 0.7800 ;
        RECT 3.9550 1.3650 4.0750 1.7250 ;
    END
    ANTENNADIFFAREA 0.1724 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.3100 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.4500 0.8750 1.5500 ;
        RECT 0.2600 1.5500 0.3700 1.6650 ;
        RECT 0.7750 1.0050 0.8750 1.4500 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5700 1.2350 0.6600 ;
      RECT 1.1450 0.6600 1.2350 0.9000 ;
      RECT 0.0700 1.8150 0.2100 1.9850 ;
      RECT 0.0700 0.9200 0.1600 1.8150 ;
      RECT 0.0700 0.6850 0.1800 0.8300 ;
      RECT 0.0700 0.8300 0.7250 0.9200 ;
      RECT 0.6350 0.6600 0.7250 0.8300 ;
      RECT 0.8400 1.7650 1.7150 1.7700 ;
      RECT 1.4150 1.7700 1.7150 1.8550 ;
      RECT 0.8400 1.6800 1.5050 1.7650 ;
      RECT 0.9650 1.0100 1.5700 1.1000 ;
      RECT 1.4800 0.4300 1.5700 1.0100 ;
      RECT 0.9650 1.1000 1.0550 1.6800 ;
      RECT 0.9650 0.8500 1.0550 1.0100 ;
      RECT 0.8550 0.7500 1.0550 0.8500 ;
      RECT 0.8400 1.7700 0.9300 1.9900 ;
      RECT 1.8400 1.2650 2.6100 1.3650 ;
      RECT 2.5100 1.3650 2.6100 1.4750 ;
      RECT 1.8400 1.3650 1.9300 1.9350 ;
      RECT 1.8400 0.6800 1.9300 1.2650 ;
      RECT 2.6300 1.5950 2.8200 1.6950 ;
      RECT 2.7300 1.1750 2.8200 1.5950 ;
      RECT 2.1250 1.0850 2.8200 1.1750 ;
      RECT 2.7300 0.8500 2.8200 1.0850 ;
      RECT 2.6700 0.6800 2.8200 0.8500 ;
      RECT 2.9200 1.6050 3.6200 1.7050 ;
      RECT 3.5200 1.1850 3.6200 1.6050 ;
      RECT 2.9200 0.6800 3.0200 1.6050 ;
      RECT 3.7300 1.0750 3.9600 1.1550 ;
      RECT 3.2950 0.9850 3.9600 1.0750 ;
      RECT 3.7300 1.1550 3.8300 1.7400 ;
      RECT 3.2950 1.0750 3.3850 1.1800 ;
      RECT 3.7850 0.6800 3.8850 0.9850 ;
      RECT 2.0200 1.8300 4.9400 1.9200 ;
      RECT 4.8500 0.9750 4.9400 1.8300 ;
      RECT 4.3500 0.8850 4.9400 0.9750 ;
      RECT 4.3500 0.6800 4.4400 0.8850 ;
      RECT 2.0200 1.4750 2.1100 1.8300 ;
      RECT 4.5300 0.6850 5.1200 0.7750 ;
      RECT 5.0300 0.7750 5.1200 1.9500 ;
      RECT 2.0500 0.5700 2.1400 0.9050 ;
      RECT 1.6600 0.4800 2.1400 0.5700 ;
      RECT 1.6600 0.5700 1.7500 1.6050 ;
      RECT 2.0500 0.9050 2.5800 0.9950 ;
      RECT 2.4900 0.5700 2.5800 0.9050 ;
      RECT 2.4900 0.4800 3.2050 0.5700 ;
      RECT 3.1150 0.5700 3.2050 0.7850 ;
      RECT 3.1150 0.8750 3.2050 1.4900 ;
      RECT 3.6050 0.4800 4.6200 0.5700 ;
      RECT 4.5300 0.5700 4.6200 0.6850 ;
      RECT 3.1150 0.7850 3.6950 0.8750 ;
      RECT 3.6050 0.5700 3.6950 0.7850 ;
  END
END SDFFQ_X0P5M_A12TH

MACRO SDFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7250 ;
        RECT 2.2800 0.3200 2.3800 0.8500 ;
        RECT 3.2150 0.3200 3.5850 0.3800 ;
        RECT 4.7400 0.3200 4.8500 0.6400 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0200 0.7250 4.1500 1.7100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.0100 5.0350 1.1900 ;
        RECT 4.9300 1.1900 5.0350 1.4450 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.2000 ;
        RECT 0.4500 1.2000 0.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 3.2600 2.0200 3.6300 2.0800 ;
        RECT 2.3150 1.9050 2.4850 2.0800 ;
        RECT 1.0700 1.8200 1.1800 2.0800 ;
        RECT 0.3350 1.6900 0.4450 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1750 1.2500 1.5350 1.3700 ;
    END
    ANTENNAGATEAREA 0.0606 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.8750 1.5500 ;
        RECT 0.7750 1.0400 0.8750 1.4500 ;
    END
    ANTENNAGATEAREA 0.0621 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5550 1.2350 0.6450 ;
      RECT 1.1450 0.6450 1.2350 0.9200 ;
      RECT 0.0450 0.8150 0.7250 0.9050 ;
      RECT 0.6350 0.6450 0.7250 0.8150 ;
      RECT 0.0450 1.6950 0.1950 1.8800 ;
      RECT 0.0450 0.9050 0.1350 1.6950 ;
      RECT 1.2700 1.8750 1.6700 1.9650 ;
      RECT 1.2700 1.7300 1.3600 1.8750 ;
      RECT 0.8300 1.6400 1.3600 1.7300 ;
      RECT 0.9650 1.0300 1.5700 1.1200 ;
      RECT 1.4800 0.4300 1.5700 1.0300 ;
      RECT 0.8300 1.7300 0.9300 1.8800 ;
      RECT 0.9650 1.1200 1.0550 1.6400 ;
      RECT 0.9650 0.9100 1.0550 1.0300 ;
      RECT 0.8550 0.8100 1.0550 0.9100 ;
      RECT 1.8400 1.1400 2.5400 1.2400 ;
      RECT 1.7600 1.8700 1.9300 1.9700 ;
      RECT 1.8400 1.2400 1.9300 1.8700 ;
      RECT 1.8400 0.6800 1.9300 1.1400 ;
      RECT 2.2000 1.5400 2.7450 1.6350 ;
      RECT 2.2000 1.3350 2.2950 1.5400 ;
      RECT 2.6500 0.7700 2.7450 1.5400 ;
      RECT 2.8750 1.6500 3.6800 1.7400 ;
      RECT 3.5900 1.0850 3.6800 1.6500 ;
      RECT 2.8750 0.9200 2.9700 1.6500 ;
      RECT 2.8750 0.7250 3.0050 0.9200 ;
      RECT 3.7700 1.5500 3.9300 1.7400 ;
      RECT 3.8400 0.7500 3.9300 1.5500 ;
      RECT 3.3050 0.6600 3.9300 0.7500 ;
      RECT 3.3050 0.7500 3.3950 1.2650 ;
      RECT 4.4300 1.6500 4.6350 1.7400 ;
      RECT 4.4300 0.5950 4.5200 1.6500 ;
      RECT 4.4300 0.5700 4.6300 0.5950 ;
      RECT 2.4700 0.4800 4.6300 0.5700 ;
      RECT 2.4700 0.5700 2.5600 0.9600 ;
      RECT 3.0950 0.5700 3.1850 1.3700 ;
      RECT 2.6850 0.4200 2.8550 0.4800 ;
      RECT 2.0400 0.9600 2.5600 1.0500 ;
      RECT 3.0600 1.3700 3.1850 1.5400 ;
      RECT 2.0400 0.5700 2.1300 0.9600 ;
      RECT 1.6600 0.4800 2.1300 0.5700 ;
      RECT 1.6600 0.5700 1.7500 1.5750 ;
      RECT 2.5950 1.8300 5.1250 1.9200 ;
      RECT 4.7450 1.8200 5.1250 1.8300 ;
      RECT 5.0250 1.6500 5.1250 1.8200 ;
      RECT 4.6400 0.8200 5.1250 0.9100 ;
      RECT 5.0250 0.4150 5.1250 0.8200 ;
      RECT 4.7450 1.5400 4.8350 1.8200 ;
      RECT 4.6400 1.4500 4.8350 1.5400 ;
      RECT 2.0200 1.6100 2.1100 1.7250 ;
      RECT 4.6400 0.9100 4.7300 1.4500 ;
      RECT 2.7300 1.9200 2.9000 1.9900 ;
      RECT 2.5950 1.8150 2.6850 1.8300 ;
      RECT 2.0200 1.7250 2.6850 1.8150 ;
  END
END SDFFQ_X1M_A12TH

MACRO SDFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6950 ;
        RECT 3.4000 0.3200 3.6100 0.3800 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9900 0.3500 1.4000 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 1.0050 5.3500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1000 1.2500 4.7250 1.3500 ;
        RECT 4.1000 1.3500 4.2000 1.7150 ;
        RECT 4.6250 1.3500 4.7250 1.7050 ;
        RECT 4.6250 0.7800 4.7250 1.2500 ;
        RECT 4.0000 0.6800 4.7250 0.7800 ;
    END
    ANTENNADIFFAREA 0.52 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5900 1.4200 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.9400 2.0550 1.1100 2.0800 ;
        RECT 2.3750 2.0300 2.5900 2.0800 ;
        RECT 0.3300 1.7350 0.4400 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1350 1.2300 1.5450 1.3500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.0500 0.7950 0.8150 0.8850 ;
      RECT 0.7250 0.8850 0.8150 1.4450 ;
      RECT 0.0500 1.7000 0.2000 1.8950 ;
      RECT 0.0500 0.8850 0.1400 1.7000 ;
      RECT 0.0500 0.5050 0.1800 0.7950 ;
      RECT 0.7700 1.7750 1.6400 1.8650 ;
      RECT 0.9350 0.8100 1.5850 0.9000 ;
      RECT 1.4950 0.4800 1.5850 0.8100 ;
      RECT 0.9350 0.9000 1.0250 1.7750 ;
      RECT 0.9350 0.6400 1.0250 0.8100 ;
      RECT 0.7600 0.5400 1.0250 0.6400 ;
      RECT 1.7300 1.8700 1.9450 1.9700 ;
      RECT 1.8550 1.2550 1.9450 1.8700 ;
      RECT 1.8550 1.1550 2.5300 1.2550 ;
      RECT 1.8550 0.7300 1.9450 1.1550 ;
      RECT 2.7200 1.5250 2.8200 1.7400 ;
      RECT 2.1500 1.4250 2.8200 1.5250 ;
      RECT 2.6300 1.3700 2.8200 1.4250 ;
      RECT 2.6300 0.6600 2.7300 1.3700 ;
      RECT 2.9400 1.6500 3.7050 1.7400 ;
      RECT 3.6150 1.0350 3.7050 1.6500 ;
      RECT 2.9400 0.6800 3.0350 1.6500 ;
      RECT 3.8000 1.0300 4.5350 1.1400 ;
      RECT 3.8550 1.1400 3.9450 1.7200 ;
      RECT 3.8000 0.9250 3.8900 1.0300 ;
      RECT 3.3700 0.8350 3.8900 0.9250 ;
      RECT 3.3700 0.9250 3.4600 1.1800 ;
      RECT 3.8000 0.6600 3.8900 0.8350 ;
      RECT 4.8200 1.5850 5.0300 1.6850 ;
      RECT 4.8200 0.5700 4.9100 1.5850 ;
      RECT 1.6750 0.4800 4.9100 0.5700 ;
      RECT 1.6750 0.5700 1.7650 1.4550 ;
      RECT 3.1500 0.5700 3.2400 1.4400 ;
      RECT 2.7800 0.4100 2.9500 0.4800 ;
      RECT 1.5750 1.4550 1.7650 1.5550 ;
      RECT 3.1500 1.4400 3.3250 1.5300 ;
      RECT 2.0350 1.8300 5.3700 1.9200 ;
      RECT 5.2800 1.6800 5.3700 1.8300 ;
      RECT 5.2800 1.5900 5.5550 1.6800 ;
      RECT 5.4650 0.5900 5.5550 1.5900 ;
      RECT 5.0000 0.5000 5.5550 0.5900 ;
      RECT 5.0000 0.5900 5.0900 1.2250 ;
      RECT 2.8350 1.9200 3.0050 1.9900 ;
      RECT 2.0350 1.6700 2.1250 1.8300 ;
  END
END SDFFQ_X2M_A12TH

MACRO SDFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4300 ;
        RECT 0.9100 0.3200 1.0100 0.6050 ;
        RECT 3.3150 0.3200 3.5250 0.3950 ;
        RECT 5.2950 0.3200 5.4150 0.6000 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1950 0.9500 1.3900 ;
        RECT 0.7700 1.0150 0.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2200 1.2900 4.8400 1.3900 ;
        RECT 4.2200 1.3900 4.3200 1.6950 ;
        RECT 4.7400 1.3900 4.8400 1.7000 ;
        RECT 4.6500 0.9250 4.7500 1.2900 ;
        RECT 4.1650 0.8250 4.8850 0.9250 ;
    END
    ANTENNADIFFAREA 0.6048 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 1.0200 5.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0600 1.3950 1.3900 ;
    END
    ANTENNAGATEAREA 0.093 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0150 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4850 0.4200 0.8000 0.5200 ;
      RECT 0.0500 1.8200 0.7650 1.9200 ;
      RECT 0.0500 0.5200 0.5850 0.6200 ;
      RECT 0.0500 0.6200 0.1500 1.8200 ;
      RECT 1.3350 1.7300 1.5050 1.9600 ;
      RECT 0.4400 1.6400 1.5050 1.7300 ;
      RECT 0.3700 0.8100 1.4700 0.9100 ;
      RECT 1.3700 0.4650 1.4700 0.8100 ;
      RECT 0.4400 0.9100 0.5300 1.6400 ;
      RECT 1.6450 1.6350 1.9100 1.7250 ;
      RECT 1.8200 0.9800 1.9100 1.6350 ;
      RECT 1.7400 0.8800 1.9100 0.9800 ;
      RECT 1.7400 0.7900 2.4500 0.8800 ;
      RECT 2.3600 0.8800 2.4500 1.2400 ;
      RECT 2.0650 1.6150 2.6300 1.7050 ;
      RECT 2.0650 1.1400 2.1550 1.6150 ;
      RECT 2.5400 0.7300 2.6300 1.6150 ;
      RECT 2.7900 0.9250 2.8900 1.6400 ;
      RECT 2.7900 0.8250 3.6050 0.9250 ;
      RECT 3.5050 0.9250 3.6050 1.2300 ;
      RECT 3.6950 1.0800 4.5550 1.1800 ;
      RECT 3.6950 1.4450 3.7950 1.7050 ;
      RECT 3.2750 1.3450 3.7950 1.4450 ;
      RECT 3.6950 1.1800 3.7950 1.3450 ;
      RECT 3.2750 1.0350 3.3750 1.3450 ;
      RECT 3.6950 0.7650 3.7950 1.0800 ;
      RECT 1.5600 0.4850 5.0850 0.5750 ;
      RECT 4.9950 0.5750 5.0850 1.7300 ;
      RECT 1.5600 1.4150 1.7300 1.5150 ;
      RECT 1.5600 0.5750 1.6500 1.4150 ;
      RECT 2.9500 0.4100 3.1200 0.4850 ;
      RECT 1.8000 1.8200 5.7550 1.9100 ;
      RECT 5.6650 0.7900 5.7550 1.8200 ;
      RECT 5.1900 0.7000 5.7550 0.7900 ;
      RECT 5.1900 0.7900 5.2800 1.2400 ;
      RECT 1.8000 1.9100 1.9200 1.9900 ;
      RECT 2.9800 1.9100 3.2200 1.9900 ;
      RECT 2.9800 1.1350 3.0700 1.8200 ;
      RECT 2.9800 1.0350 3.1600 1.1350 ;
  END
END SDFFQ_X3M_A12TH

MACRO SDFFQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4300 ;
        RECT 0.9100 0.3200 1.0100 0.5800 ;
        RECT 3.3350 0.3200 3.5450 0.3850 ;
        RECT 5.6950 0.3200 5.7950 0.7050 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1950 0.9500 1.3900 ;
        RECT 0.7700 1.0100 0.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.8600 4.9800 1.2900 ;
        RECT 4.3600 1.2900 4.9800 1.3900 ;
        RECT 4.3050 0.7600 4.9800 0.8600 ;
        RECT 4.3600 1.3900 4.4600 1.7000 ;
        RECT 4.8800 1.3900 4.9800 1.7000 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8450 1.0200 5.9650 1.5000 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0600 1.3950 1.3900 ;
    END
    ANTENNAGATEAREA 0.0945 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0150 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0795 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3950 0.4150 0.7750 0.5150 ;
      RECT 0.0500 1.8200 0.7650 1.9200 ;
      RECT 0.0500 0.5700 0.4950 0.6700 ;
      RECT 0.3950 0.5150 0.4950 0.5700 ;
      RECT 0.0500 0.6700 0.1500 1.8200 ;
      RECT 1.3350 1.7300 1.5050 1.9650 ;
      RECT 0.4400 1.6400 1.5050 1.7300 ;
      RECT 0.3700 0.8050 1.4700 0.9050 ;
      RECT 1.3700 0.4550 1.4700 0.8050 ;
      RECT 0.4400 0.9050 0.5300 1.6400 ;
      RECT 1.6500 1.5300 1.9100 1.6200 ;
      RECT 1.8200 0.8750 1.9100 1.5300 ;
      RECT 1.7400 0.7750 1.9100 0.8750 ;
      RECT 1.7400 0.6850 2.4400 0.7750 ;
      RECT 2.3500 0.7750 2.4400 1.2400 ;
      RECT 2.0650 1.5450 2.6200 1.6350 ;
      RECT 2.0650 1.0200 2.1550 1.5450 ;
      RECT 2.5300 0.7300 2.6200 1.5450 ;
      RECT 2.7200 0.9300 2.8200 1.7050 ;
      RECT 2.7200 0.8300 3.6500 0.9300 ;
      RECT 3.5500 0.9300 3.6500 1.4700 ;
      RECT 3.7400 1.0800 4.7300 1.1800 ;
      RECT 3.2950 1.6100 3.8400 1.7100 ;
      RECT 3.7400 1.1800 3.8400 1.6100 ;
      RECT 3.2950 1.0500 3.3950 1.6100 ;
      RECT 3.7400 0.7300 3.8400 1.0800 ;
      RECT 1.5600 0.4850 5.4850 0.5750 ;
      RECT 5.3950 0.5750 5.4850 1.7200 ;
      RECT 1.5600 1.3050 1.7300 1.4050 ;
      RECT 1.5600 0.5750 1.6500 1.3050 ;
      RECT 3.0250 0.4100 3.1950 0.4850 ;
      RECT 1.8000 1.8150 6.1550 1.9050 ;
      RECT 6.0650 0.9050 6.1550 1.8150 ;
      RECT 5.5800 0.8150 6.1550 0.9050 ;
      RECT 6.0250 0.5200 6.1550 0.8150 ;
      RECT 5.5800 0.9050 5.6700 1.4600 ;
      RECT 1.8000 1.9050 1.9200 1.9900 ;
      RECT 3.2300 1.9050 3.3750 1.9900 ;
      RECT 3.0650 1.0350 3.1650 1.8150 ;
  END
END SDFFQ_X4M_A12TH

MACRO PREICG_X0P6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 2.6700 0.3200 2.7600 0.6900 ;
        RECT 0.3800 0.3200 0.4700 0.6150 ;
        RECT 1.2450 0.3200 1.3350 0.5250 ;
        RECT 3.2300 0.3200 3.3200 0.8350 ;
        RECT 2.6700 0.6900 2.8400 0.7800 ;
        RECT 0.3000 0.6150 0.4700 0.7050 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8800 0.1500 1.6200 ;
        RECT 0.0600 1.6200 0.1850 1.7100 ;
        RECT 0.0600 0.7100 0.1700 0.8800 ;
        RECT 0.0950 1.7100 0.1850 1.9900 ;
    END
    ANTENNADIFFAREA 0.138575 ;
  END ECK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7800 1.0500 3.2150 1.1500 ;
        RECT 3.1250 1.1500 3.2150 1.2300 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7450 1.2500 1.0400 1.3700 ;
        RECT 0.9500 1.3700 1.0400 1.4350 ;
        RECT 0.9500 1.4350 1.5650 1.5250 ;
        RECT 1.4750 1.5250 1.5650 1.7650 ;
        RECT 1.4750 1.7650 1.9000 1.8550 ;
        RECT 1.8100 1.8550 1.9000 1.8800 ;
        RECT 1.8100 1.8800 2.2250 1.9700 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.4100 3.1600 1.5100 ;
        RECT 2.8500 1.5100 2.9500 1.5900 ;
        RECT 2.8500 1.2650 2.9400 1.4100 ;
    END
    ANTENNAGATEAREA 0.0372 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.9400 1.9000 1.0300 2.0800 ;
        RECT 2.5800 1.8800 2.7500 2.0800 ;
        RECT 0.3550 1.8450 0.4450 2.0800 ;
        RECT 1.2150 1.6150 1.3850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.7950 0.9550 0.8850 ;
      RECT 0.8650 0.7100 0.9550 0.7950 ;
      RECT 0.5550 1.7550 0.6450 1.8450 ;
      RECT 0.3400 1.6650 0.6450 1.7550 ;
      RECT 0.3400 1.5450 0.4300 1.6650 ;
      RECT 0.2750 1.3750 0.4300 1.5450 ;
      RECT 0.3400 0.8850 0.4300 1.3750 ;
      RECT 0.5550 1.8450 0.8300 1.9350 ;
      RECT 0.5200 0.9750 1.4100 1.0650 ;
      RECT 1.3200 0.8850 1.4100 0.9750 ;
      RECT 0.7500 1.6150 1.0950 1.7050 ;
      RECT 1.0450 0.5000 1.1350 0.9750 ;
      RECT 0.9450 0.4100 1.1350 0.5000 ;
      RECT 0.5200 1.0650 0.6100 1.4850 ;
      RECT 0.7500 1.5750 0.8400 1.6150 ;
      RECT 0.5200 1.4850 0.8400 1.5750 ;
      RECT 1.6900 1.5850 1.8600 1.6750 ;
      RECT 1.6900 1.3450 1.7800 1.5850 ;
      RECT 1.1400 1.2550 1.7800 1.3450 ;
      RECT 1.5000 0.9850 1.5900 1.2550 ;
      RECT 1.5000 0.8950 1.7400 0.9850 ;
      RECT 1.6500 0.5000 1.7400 0.8950 ;
      RECT 1.6500 0.4100 1.8750 0.5000 ;
      RECT 1.1400 1.1750 1.2300 1.2550 ;
      RECT 2.2450 1.5200 2.4150 1.6100 ;
      RECT 2.2450 1.1650 2.3350 1.5200 ;
      RECT 1.7000 1.0900 2.3350 1.1650 ;
      RECT 1.7000 1.0750 2.3750 1.0900 ;
      RECT 2.1500 0.9900 2.3750 1.0750 ;
      RECT 2.2850 0.7350 2.3750 0.9900 ;
      RECT 1.9900 1.7000 3.3200 1.7700 ;
      RECT 2.5250 1.6800 3.3200 1.7000 ;
      RECT 3.2300 1.6000 3.3200 1.6800 ;
      RECT 1.9900 1.7700 2.6150 1.7900 ;
      RECT 1.9900 1.6150 2.0800 1.7000 ;
      RECT 2.5250 0.9600 2.6150 1.6800 ;
      RECT 2.4750 0.5700 2.5650 0.8700 ;
      RECT 1.9900 0.4800 2.5650 0.5700 ;
      RECT 1.9900 0.4250 2.1600 0.4800 ;
      RECT 2.4750 0.8700 3.0600 0.9600 ;
      RECT 2.9700 0.7350 3.0600 0.8700 ;
  END
END PREICG_X0P6B_A12TH

MACRO PREICG_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9000 ;
        RECT 1.3250 0.3200 1.4150 0.5850 ;
        RECT 2.5800 0.3200 2.7500 0.5200 ;
        RECT 3.1750 0.3200 3.3550 0.7500 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1900 1.0500 2.6050 1.1600 ;
        RECT 2.5150 1.1600 2.6050 1.5600 ;
        RECT 2.1550 1.5600 2.6050 1.6500 ;
        RECT 2.1550 1.6500 2.2450 1.8300 ;
        RECT 0.8800 1.8300 2.2450 1.9200 ;
        RECT 0.8800 1.7550 0.9700 1.8300 ;
        RECT 0.8150 1.6650 0.9700 1.7550 ;
        RECT 0.8150 1.5450 0.9050 1.6650 ;
    END
    ANTENNAGATEAREA 0.0735 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.1500 1.5350 ;
        RECT 0.0600 1.5350 0.1700 1.6250 ;
        RECT 0.0600 0.9100 0.1700 1.0000 ;
        RECT 0.0800 1.6250 0.1700 1.9050 ;
        RECT 0.0800 0.7900 0.1700 0.9100 ;
    END
    ANTENNADIFFAREA 0.1528 ;
  END ECK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7850 1.2500 3.1550 1.3500 ;
        RECT 3.0550 1.0200 3.1550 1.2500 ;
    END
    ANTENNAGATEAREA 0.0297 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5600 0.8500 2.8800 0.9500 ;
        RECT 2.7800 0.9500 2.8800 1.1400 ;
    END
    ANTENNAGATEAREA 0.0381 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.9300 2.0100 1.1400 2.0800 ;
        RECT 0.3400 1.8250 0.4300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3050 0.9900 1.0100 1.0800 ;
      RECT 0.9200 0.7800 1.0100 0.9900 ;
      RECT 0.6000 1.8700 0.7900 1.9600 ;
      RECT 0.6000 1.5550 0.6900 1.8700 ;
      RECT 0.3050 1.4650 0.6900 1.5550 ;
      RECT 0.3050 1.4450 0.3950 1.4650 ;
      RECT 0.2400 1.2350 0.3950 1.4450 ;
      RECT 0.3050 1.0800 0.3950 1.2350 ;
      RECT 1.0800 1.4700 1.6750 1.5600 ;
      RECT 1.0800 1.6500 1.2700 1.7400 ;
      RECT 1.0800 1.5600 1.1900 1.6500 ;
      RECT 1.0800 1.3750 1.1900 1.4700 ;
      RECT 0.5550 1.2850 1.1900 1.3750 ;
      RECT 1.1000 0.6000 1.1900 1.2850 ;
      RECT 1.0200 0.5100 1.1900 0.6000 ;
      RECT 1.0200 0.4100 1.1100 0.5100 ;
      RECT 0.5550 1.1700 0.6450 1.2850 ;
      RECT 1.7650 1.6500 2.0450 1.7400 ;
      RECT 1.7650 1.3600 1.8550 1.6500 ;
      RECT 1.2800 1.2700 1.8550 1.3600 ;
      RECT 1.2800 1.1500 1.3700 1.2700 ;
      RECT 1.5250 0.5900 1.6150 1.2700 ;
      RECT 1.5250 0.5000 1.9900 0.5900 ;
      RECT 1.9000 0.4100 1.9900 0.5000 ;
      RECT 2.3350 1.3600 2.4250 1.4500 ;
      RECT 1.9450 1.2700 2.4250 1.3600 ;
      RECT 1.9450 0.7700 2.2750 0.8600 ;
      RECT 1.8950 0.6800 2.2750 0.7700 ;
      RECT 2.1850 0.6500 2.2750 0.6800 ;
      RECT 1.9450 1.1800 2.0350 1.2700 ;
      RECT 1.7250 1.0900 2.0350 1.1800 ;
      RECT 1.9450 0.8600 2.0350 1.0900 ;
      RECT 2.3550 1.7400 3.3550 1.8300 ;
      RECT 3.2650 1.5300 3.3550 1.7400 ;
      RECT 3.1550 1.4400 3.3550 1.5300 ;
      RECT 3.2650 0.9300 3.3550 1.4400 ;
      RECT 2.9950 0.8400 3.3550 0.9300 ;
      RECT 2.3650 0.5400 2.4550 0.6200 ;
      RECT 2.1000 0.4500 2.4550 0.5400 ;
      RECT 2.9950 0.7600 3.0850 0.8400 ;
      RECT 2.8450 0.7100 3.0850 0.7600 ;
      RECT 2.3650 0.6200 3.0850 0.7100 ;
  END
END PREICG_X0P7B_A12TH

MACRO PREICG_X0P8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.9800 ;
        RECT 1.3750 0.3200 1.4650 0.6000 ;
        RECT 2.5800 0.3200 2.7500 0.4550 ;
        RECT 3.1650 0.3200 3.3550 0.7300 ;
    END
  END VSS

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 1.2100 3.1500 1.4100 ;
        RECT 3.0500 1.0000 3.1650 1.2100 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.2700 2.9500 1.5900 ;
        RECT 2.8050 1.1900 2.9500 1.2700 ;
        RECT 2.8050 1.0200 2.8950 1.1900 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END SE

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9800 0.1500 1.4450 ;
        RECT 0.0600 1.4450 0.1700 1.5350 ;
        RECT 0.0600 0.8900 0.1700 0.9800 ;
        RECT 0.0800 1.5350 0.1700 1.8150 ;
        RECT 0.0800 0.6100 0.1700 0.8900 ;
    END
    ANTENNADIFFAREA 0.1736 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.9300 2.0000 1.1400 2.0800 ;
        RECT 0.3400 1.8200 0.4300 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0850 1.0500 2.6350 1.1500 ;
        RECT 2.5350 1.1500 2.6350 1.5450 ;
        RECT 2.1050 1.5450 2.6350 1.6350 ;
        RECT 2.1050 1.6350 2.1950 1.8200 ;
        RECT 0.8800 1.8200 2.1950 1.9100 ;
        RECT 0.8800 1.7100 0.9700 1.8200 ;
        RECT 0.7750 1.6200 0.9700 1.7100 ;
        RECT 0.7750 1.5000 0.8650 1.6200 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.2800 1.0700 0.9700 1.1600 ;
      RECT 0.8800 0.7900 0.9700 1.0700 ;
      RECT 0.5600 1.6400 0.6500 1.8350 ;
      RECT 0.2800 1.5500 0.6500 1.6400 ;
      RECT 0.2800 1.1600 0.3700 1.5500 ;
      RECT 0.5600 1.8350 0.7900 1.9250 ;
      RECT 1.0800 1.3400 1.5900 1.3500 ;
      RECT 0.5350 1.2600 1.5900 1.3400 ;
      RECT 1.5000 1.1400 1.5900 1.2600 ;
      RECT 1.0800 1.3500 1.1700 1.6800 ;
      RECT 0.5350 1.2500 1.1500 1.2600 ;
      RECT 1.0600 0.5550 1.1500 1.2500 ;
      RECT 0.9950 0.4650 1.2050 0.5550 ;
      RECT 0.5350 1.3400 0.6250 1.4600 ;
      RECT 1.8050 1.6400 1.9950 1.7300 ;
      RECT 1.7000 1.5500 1.8950 1.6400 ;
      RECT 1.7000 1.0500 1.7900 1.5500 ;
      RECT 1.2650 0.9600 1.7900 1.0500 ;
      RECT 1.7000 0.5550 1.7900 0.9600 ;
      RECT 1.7000 0.4650 2.0450 0.5550 ;
      RECT 1.2650 0.8400 1.3550 0.9600 ;
      RECT 1.9000 1.2600 2.4450 1.3500 ;
      RECT 2.3550 1.3500 2.4450 1.4350 ;
      RECT 1.9000 0.8150 2.1700 0.9050 ;
      RECT 2.0100 0.7250 2.4250 0.8150 ;
      RECT 1.9000 1.3500 1.9900 1.4600 ;
      RECT 1.9000 0.9050 1.9900 1.2600 ;
      RECT 2.3050 1.7250 3.3200 1.8150 ;
      RECT 3.2300 1.6100 3.3200 1.7250 ;
      RECT 3.2300 1.5200 3.3500 1.6100 ;
      RECT 3.2600 0.9100 3.3500 1.5200 ;
      RECT 2.9650 0.8200 3.3500 0.9100 ;
      RECT 2.9650 0.6350 3.0550 0.8200 ;
      RECT 2.3750 0.5550 3.0550 0.6350 ;
      RECT 2.1600 0.5450 3.0550 0.5550 ;
      RECT 2.1600 0.4650 2.4650 0.5450 ;
  END
END PREICG_X0P8B_A12TH

MACRO PREICG_X11B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7400 ;
        RECT 0.8600 0.3200 0.9600 0.7400 ;
        RECT 1.8050 0.3200 2.1750 0.3400 ;
        RECT 3.7900 0.3200 3.8900 0.6300 ;
        RECT 4.7500 0.3200 4.8500 0.6300 ;
        RECT 5.3450 0.3200 5.4450 0.5900 ;
        RECT 5.8650 0.3200 5.9650 0.5900 ;
        RECT 6.3850 0.3200 6.4850 0.5900 ;
        RECT 6.9050 0.3200 7.0050 0.5900 ;
        RECT 7.4250 0.3200 7.5250 0.5900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 4.8250 1.7700 4.9250 2.0800 ;
        RECT 5.3450 1.7700 5.4450 2.0800 ;
        RECT 5.8650 1.7700 5.9650 2.0800 ;
        RECT 6.3850 1.7700 6.4850 2.0800 ;
        RECT 6.9050 1.7700 7.0050 2.0800 ;
        RECT 7.4250 1.7700 7.5250 2.0800 ;
        RECT 3.3300 1.7450 3.4300 2.0800 ;
        RECT 4.0300 1.7450 4.1300 2.0800 ;
        RECT 4.5500 1.7450 4.6500 2.0800 ;
        RECT 2.0600 1.7100 2.1600 2.0800 ;
        RECT 2.8050 1.5250 2.9050 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1200 1.0500 4.5750 1.1500 ;
        RECT 3.1200 0.5800 3.2200 1.0500 ;
        RECT 1.3150 0.4800 3.2200 0.5800 ;
        RECT 1.3150 0.5800 1.4150 1.4350 ;
        RECT 1.5600 0.4600 1.7300 0.4800 ;
    END
    ANTENNAGATEAREA 0.4407 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2200 0.8450 7.3800 1.2200 ;
        RECT 5.0850 1.2200 7.3800 1.3800 ;
        RECT 5.0850 0.6850 7.3800 0.8450 ;
        RECT 5.0850 1.3800 5.1850 1.7200 ;
        RECT 5.6050 1.3800 5.7050 1.7200 ;
        RECT 6.1250 1.3800 6.2250 1.7200 ;
        RECT 6.6450 1.3800 6.7450 1.7200 ;
        RECT 7.1650 1.3800 7.2650 1.7200 ;
        RECT 5.0900 0.4900 5.1800 0.6850 ;
        RECT 5.6100 0.4900 5.7000 0.6850 ;
        RECT 6.1300 0.4900 6.2200 0.6850 ;
        RECT 6.6500 0.4900 6.7400 0.6850 ;
        RECT 7.1700 0.4900 7.2600 0.6850 ;
    END
    ANTENNADIFFAREA 1.62295 ;
  END ECK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.2400 0.8150 1.3600 ;
    END
    ANTENNAGATEAREA 0.1368 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 1.0500 1.0250 1.1500 ;
        RECT 0.9250 1.1500 1.0250 1.2500 ;
    END
    ANTENNAGATEAREA 0.1068 ;
  END E
  OBS
    LAYER M1 ;
      RECT 0.2850 1.6500 1.0050 1.7400 ;
      RECT 0.0750 1.8300 1.2250 1.9200 ;
      RECT 1.1350 0.9400 1.2250 1.8300 ;
      RECT 0.0750 0.8500 1.2250 0.9400 ;
      RECT 1.1350 0.5650 1.2250 0.8500 ;
      RECT 0.0750 1.7100 0.1750 1.8300 ;
      RECT 0.0750 0.5500 0.1750 0.8500 ;
      RECT 0.5950 0.5300 0.6950 0.8500 ;
      RECT 1.3550 1.5950 1.6150 1.6850 ;
      RECT 1.5250 1.1350 1.6150 1.5950 ;
      RECT 1.5250 1.0450 2.2250 1.1350 ;
      RECT 2.1350 0.9450 2.2250 1.0450 ;
      RECT 1.5250 0.6850 1.6150 1.0450 ;
      RECT 1.7550 1.4900 2.6550 1.5800 ;
      RECT 2.5350 1.5800 2.6550 1.9450 ;
      RECT 2.5650 0.9400 2.6550 1.4900 ;
      RECT 2.5150 0.8500 2.6850 0.9400 ;
      RECT 1.5550 1.8450 1.8450 1.9350 ;
      RECT 1.7550 1.5800 1.8450 1.8450 ;
      RECT 2.9200 1.2400 4.7750 1.3300 ;
      RECT 4.6850 1.0050 4.7750 1.2400 ;
      RECT 1.8250 1.3100 2.4550 1.4000 ;
      RECT 2.3150 0.7600 2.4050 1.3100 ;
      RECT 2.2450 0.6700 3.0100 0.7600 ;
      RECT 2.9200 0.7600 3.0100 1.2400 ;
      RECT 4.8850 0.9550 6.9650 1.0550 ;
      RECT 3.0700 1.5300 3.1700 1.8800 ;
      RECT 3.5900 1.5300 3.6900 1.8800 ;
      RECT 3.3300 0.4650 3.4300 0.8100 ;
      RECT 4.2900 1.5300 4.3900 1.8800 ;
      RECT 4.2900 0.4650 4.3900 0.8100 ;
      RECT 3.0700 1.4400 4.9750 1.5300 ;
      RECT 4.8850 1.0550 4.9750 1.4400 ;
      RECT 4.8850 0.9000 4.9750 0.9550 ;
      RECT 3.3300 0.8100 4.9750 0.9000 ;
  END
END PREICG_X11B_A12TH

MACRO PREICG_X13B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 9.6450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.5800 ;
        RECT 0.8700 0.3200 0.9700 0.5800 ;
        RECT 3.0650 0.3200 3.2350 0.3750 ;
        RECT 3.6200 0.3200 3.7900 0.3400 ;
        RECT 4.6400 0.3200 4.7400 0.6650 ;
        RECT 5.5600 0.3200 5.6600 0.6650 ;
        RECT 6.2700 0.3200 6.3700 0.6650 ;
        RECT 6.7900 0.3200 6.8900 0.6000 ;
        RECT 7.3100 0.3200 7.4100 0.5450 ;
        RECT 7.8300 0.3200 7.9300 0.5450 ;
        RECT 8.3500 0.3200 8.4500 0.5450 ;
        RECT 8.8700 0.3200 8.9700 0.5550 ;
        RECT 9.3900 0.3200 9.4900 0.5550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 9.6450 2.7200 ;
        RECT 0.5750 1.8950 0.7450 2.0800 ;
        RECT 3.1000 1.7900 3.2000 2.0800 ;
        RECT 6.1250 1.7700 6.2250 2.0800 ;
        RECT 6.7900 1.7700 6.8900 2.0800 ;
        RECT 7.3100 1.7700 7.4100 2.0800 ;
        RECT 7.8300 1.7700 7.9300 2.0800 ;
        RECT 8.3500 1.7700 8.4500 2.0800 ;
        RECT 8.8700 1.7700 8.9700 2.0800 ;
        RECT 9.3900 1.7700 9.4900 2.0800 ;
        RECT 4.1450 1.7450 4.2450 2.0800 ;
        RECT 4.8400 1.7300 4.9400 2.0800 ;
        RECT 5.3600 1.7300 5.4600 2.0800 ;
        RECT 2.5250 1.6700 2.6250 2.0800 ;
    END
  END VDD

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8500 1.0400 0.9500 ;
        RECT 0.2500 0.9500 0.3500 1.1500 ;
        RECT 0.9400 0.9500 1.0400 1.2500 ;
    END
    ANTENNAGATEAREA 0.1218 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0400 0.8300 1.1600 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END SE

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2100 0.8850 9.3900 1.2500 ;
        RECT 6.5300 1.2500 9.3900 1.4300 ;
        RECT 6.5300 0.7050 9.3900 0.8850 ;
        RECT 6.5300 1.4300 6.6300 1.7200 ;
        RECT 7.0500 1.4300 7.1500 1.7200 ;
        RECT 7.5700 1.4300 7.6700 1.7200 ;
        RECT 8.0900 1.4300 8.1900 1.7200 ;
        RECT 8.6100 1.4300 8.7100 1.7200 ;
        RECT 9.1300 1.4300 9.2300 1.7200 ;
        RECT 6.5300 0.4950 6.6300 0.7050 ;
        RECT 7.0500 0.4550 7.1500 0.7050 ;
        RECT 7.5700 0.4550 7.6700 0.7050 ;
        RECT 8.0900 0.4550 8.1900 0.7050 ;
        RECT 8.6100 0.4550 8.7100 0.7050 ;
        RECT 9.1300 0.4550 9.2300 0.7050 ;
    END
    ANTENNADIFFAREA 1.92955 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9350 1.0500 6.0850 1.1500 ;
        RECT 3.9350 0.5800 4.0350 1.0500 ;
        RECT 1.8700 0.4800 4.0350 0.5800 ;
        RECT 1.8700 0.5800 1.9700 1.3450 ;
        RECT 1.6300 1.3450 1.9700 1.4450 ;
    END
    ANTENNAGATEAREA 0.5118 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 2.0600 1.0800 3.0600 1.1700 ;
      RECT 1.3900 1.5950 2.1500 1.6850 ;
      RECT 2.0600 1.1700 2.1500 1.5950 ;
      RECT 2.0600 0.7050 2.1500 1.0800 ;
      RECT 1.4300 0.6900 1.5200 1.5950 ;
      RECT 2.2550 1.4900 3.5750 1.5800 ;
      RECT 3.4850 0.9400 3.5750 1.4900 ;
      RECT 3.4050 0.8500 3.5750 0.9400 ;
      RECT 2.0750 1.8450 2.3450 1.9350 ;
      RECT 2.2550 1.5800 2.3450 1.8450 ;
      RECT 3.7350 1.2400 5.6800 1.3300 ;
      RECT 2.3150 1.3100 3.2800 1.4000 ;
      RECT 3.1900 0.7600 3.2800 1.3100 ;
      RECT 2.7850 0.6700 3.8250 0.7600 ;
      RECT 3.7350 0.7600 3.8250 1.2400 ;
      RECT 6.2800 0.9950 8.9500 1.0950 ;
      RECT 3.8850 1.5700 3.9850 1.9100 ;
      RECT 4.4050 1.5700 4.5050 1.9100 ;
      RECT 4.1450 0.4700 4.2450 0.8100 ;
      RECT 5.1000 1.5700 5.2000 1.9100 ;
      RECT 5.1000 0.4700 5.2000 0.8100 ;
      RECT 5.7600 1.5700 5.8600 1.9650 ;
      RECT 6.0200 0.4700 6.1200 0.8100 ;
      RECT 3.8850 1.4800 6.3700 1.5700 ;
      RECT 6.2800 1.0950 6.3700 1.4800 ;
      RECT 6.2800 0.9000 6.3700 0.9950 ;
      RECT 4.1450 0.8100 6.3700 0.9000 ;
      RECT 0.2950 1.5000 1.0200 1.5900 ;
      RECT 1.1500 1.8050 1.8400 1.8950 ;
      RECT 1.1500 0.4800 1.7800 0.5700 ;
      RECT 1.6900 0.5700 1.7800 0.8900 ;
      RECT 1.1500 1.7700 1.2400 1.8050 ;
      RECT 0.0500 1.6800 1.2400 1.7700 ;
      RECT 1.1500 0.7600 1.2400 1.6800 ;
      RECT 0.0550 0.6700 1.2400 0.7600 ;
      RECT 1.1500 0.5700 1.2400 0.6700 ;
      RECT 0.0550 0.4700 0.2250 0.6700 ;
      RECT 0.5750 0.4700 0.7450 0.6700 ;
  END
END PREICG_X13B_A12TH

MACRO PREICG_X16B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 10.6450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.7150 ;
        RECT 0.6100 0.3200 0.7100 0.5400 ;
        RECT 1.1450 0.3200 1.2450 0.5400 ;
        RECT 4.7300 0.3200 4.8300 0.6300 ;
        RECT 5.6500 0.3200 5.7500 0.6300 ;
        RECT 6.6000 0.3200 6.7000 0.6300 ;
    END
  END VSS

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0450 0.9000 1.1550 ;
    END
    ANTENNAGATEAREA 0.1446 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0500 6.3700 1.1500 ;
        RECT 4.0500 0.5800 4.1500 1.0500 ;
        RECT 1.9250 0.4800 4.1500 0.5800 ;
        RECT 1.9250 0.5800 2.0250 1.2900 ;
        RECT 3.4000 0.4100 3.5700 0.4800 ;
        RECT 1.9250 1.2900 2.0950 1.3800 ;
    END
    ANTENNAGATEAREA 0.6564 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.9900 0.7650 10.2100 1.2900 ;
        RECT 6.9250 1.2900 10.2100 1.4750 ;
        RECT 6.9200 0.5450 10.2100 0.7650 ;
        RECT 6.9200 1.4750 10.2100 1.5100 ;
        RECT 7.4050 0.4150 7.5750 0.5450 ;
        RECT 7.9250 0.4150 8.0950 0.5450 ;
        RECT 8.4450 0.4150 8.6150 0.5450 ;
        RECT 8.9650 0.4150 9.1350 0.5450 ;
        RECT 9.4850 0.4150 9.6550 0.5450 ;
        RECT 10.0050 0.4150 10.1750 0.5450 ;
        RECT 6.9200 1.5100 7.0200 1.9050 ;
        RECT 7.4400 1.5100 7.5400 1.7200 ;
        RECT 7.9600 1.5100 8.0600 1.7200 ;
        RECT 8.4800 1.5100 8.5800 1.7200 ;
        RECT 9.0000 1.5100 9.1000 1.7200 ;
        RECT 9.5200 1.5100 9.6200 1.7200 ;
        RECT 10.0400 1.5100 10.1400 1.8350 ;
    END
    ANTENNADIFFAREA 2.2735 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 10.6450 2.7200 ;
        RECT 1.1100 2.0100 1.2800 2.0800 ;
        RECT 5.8500 1.7700 5.9500 2.0800 ;
        RECT 6.4900 1.7700 6.5900 2.0800 ;
        RECT 7.1800 1.7700 7.2800 2.0800 ;
        RECT 7.7000 1.7700 7.8000 2.0800 ;
        RECT 8.2200 1.7700 8.3200 2.0800 ;
        RECT 8.7400 1.7700 8.8400 2.0800 ;
        RECT 9.2600 1.7700 9.3600 2.0800 ;
        RECT 9.7800 1.7700 9.8800 2.0800 ;
        RECT 10.3000 1.7700 10.4000 2.0800 ;
        RECT 0.0900 1.7550 0.1900 2.0800 ;
        RECT 4.2500 1.7150 4.3500 2.0800 ;
        RECT 4.9300 1.7150 5.0300 2.0800 ;
        RECT 5.4500 1.7150 5.5500 2.0800 ;
        RECT 2.7950 1.6700 2.8950 2.0800 ;
        RECT 3.3350 1.6700 3.4350 2.0800 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.2500 1.1700 1.3500 ;
        RECT 0.1950 1.0800 0.2950 1.2500 ;
        RECT 1.0700 1.0800 1.1700 1.2500 ;
    END
    ANTENNAGATEAREA 0.186 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.3500 1.8300 1.5400 1.9200 ;
      RECT 0.3500 1.5000 0.4500 1.8300 ;
      RECT 1.9350 1.7400 2.1050 1.9500 ;
      RECT 0.5600 1.6500 2.1050 1.7400 ;
      RECT 1.2850 0.7200 1.3750 1.6500 ;
      RECT 0.3150 0.6300 1.8350 0.7200 ;
      RECT 1.7450 0.7200 1.8350 0.8650 ;
      RECT 1.7450 0.4550 1.8350 0.6300 ;
      RECT 0.3150 0.4300 0.4850 0.6300 ;
      RECT 0.8500 0.4300 1.0200 0.6300 ;
      RECT 2.2350 1.0800 3.1700 1.1700 ;
      RECT 2.2350 1.5600 2.3250 1.7100 ;
      RECT 1.4850 1.4700 2.3250 1.5600 ;
      RECT 2.2350 1.1700 2.3250 1.4700 ;
      RECT 2.2350 0.9550 2.3250 1.0800 ;
      RECT 2.1150 0.8650 2.3250 0.9550 ;
      RECT 2.1150 0.6900 2.2050 0.8650 ;
      RECT 1.4850 0.8100 1.5750 1.4700 ;
      RECT 2.5650 1.4900 3.7000 1.5800 ;
      RECT 3.6100 1.5800 3.7000 1.7750 ;
      RECT 3.6100 0.9400 3.7000 1.4900 ;
      RECT 3.4600 0.8500 3.7000 0.9400 ;
      RECT 2.3400 1.8450 2.6550 1.9350 ;
      RECT 2.5650 1.5800 2.6550 1.8450 ;
      RECT 3.8500 1.2400 6.6000 1.3300 ;
      RECT 2.5250 1.3100 3.3500 1.4000 ;
      RECT 3.2600 0.7600 3.3500 1.3100 ;
      RECT 2.8550 0.6700 3.9400 0.7600 ;
      RECT 3.8500 0.7600 3.9400 1.2400 ;
      RECT 6.7100 0.8800 9.7500 0.9700 ;
      RECT 3.9900 1.4400 6.8000 1.5300 ;
      RECT 6.7100 0.9700 6.8000 1.4400 ;
      RECT 6.7100 0.8700 6.8000 0.8800 ;
      RECT 4.2700 0.7800 6.8000 0.8700 ;
      RECT 3.9900 1.5300 4.0900 1.8800 ;
      RECT 4.5100 1.5300 4.6100 1.8800 ;
      RECT 4.2700 0.4250 4.3700 0.7800 ;
      RECT 5.1900 1.5300 5.2900 1.8800 ;
      RECT 5.1900 0.4250 5.2900 0.7800 ;
      RECT 6.1100 1.5300 6.2100 1.9350 ;
      RECT 6.1100 0.4250 6.2100 0.7800 ;
  END
END PREICG_X16B_A12TH

MACRO PREICG_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3850 0.3200 0.4750 0.8000 ;
        RECT 1.4300 0.3200 1.5200 0.5550 ;
        RECT 3.2300 0.3200 3.3200 0.5200 ;
    END
  END VSS

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8750 0.8100 3.1650 0.9100 ;
        RECT 3.0500 0.9100 3.1650 1.0850 ;
    END
    ANTENNAGATEAREA 0.0321 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1900 1.0500 2.5950 1.1500 ;
        RECT 2.4950 1.1500 2.5950 1.5250 ;
        RECT 2.2100 1.5250 2.5950 1.6150 ;
        RECT 2.2100 1.6150 2.3000 1.8300 ;
        RECT 0.8450 1.8300 2.3000 1.9200 ;
        RECT 0.8450 1.2500 0.9350 1.8300 ;
    END
    ANTENNAGATEAREA 0.0837 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8000 0.1500 1.2800 ;
        RECT 0.0600 1.2800 0.1700 1.3700 ;
        RECT 0.0600 0.7100 0.1700 0.8000 ;
        RECT 0.0800 1.3700 0.1700 1.6500 ;
        RECT 0.0800 0.4300 0.1700 0.7100 ;
    END
    ANTENNADIFFAREA 0.2184 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.9400 2.0100 1.1500 2.0800 ;
        RECT 0.3400 1.8550 0.4300 2.0800 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8100 1.0200 2.9500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 0.2400 0.8900 0.9700 0.9800 ;
      RECT 0.8800 0.6100 0.9700 0.8900 ;
      RECT 0.6650 1.4600 0.7550 1.6850 ;
      RECT 0.2600 1.3700 0.7550 1.4600 ;
      RECT 0.2600 1.1000 0.3500 1.3700 ;
      RECT 0.2400 0.9800 0.3500 1.1000 ;
      RECT 1.0800 0.9300 1.6000 1.0200 ;
      RECT 1.5100 1.0200 1.6000 1.1150 ;
      RECT 1.0800 1.6450 1.3450 1.7350 ;
      RECT 1.0800 1.1600 1.1700 1.6450 ;
      RECT 0.5350 1.0700 1.1700 1.1600 ;
      RECT 1.0800 1.0200 1.1700 1.0700 ;
      RECT 1.0800 0.5200 1.1700 0.9300 ;
      RECT 1.0800 0.4300 1.2950 0.5200 ;
      RECT 0.5350 1.1600 0.6250 1.2800 ;
      RECT 1.6900 1.6300 2.1200 1.7200 ;
      RECT 1.6900 1.4050 1.7800 1.6300 ;
      RECT 1.2600 1.3150 1.7800 1.4050 ;
      RECT 1.6900 0.6700 1.7800 1.3150 ;
      RECT 1.6900 0.5800 1.9500 0.6700 ;
      RECT 1.8600 0.5200 1.9500 0.5800 ;
      RECT 1.8600 0.4300 2.1000 0.5200 ;
      RECT 1.8900 1.3250 2.4050 1.4150 ;
      RECT 1.8900 0.7800 2.2600 0.8700 ;
      RECT 2.1700 0.6900 2.4250 0.7800 ;
      RECT 1.8900 0.8700 1.9800 1.3250 ;
      RECT 2.3900 1.7250 3.3200 1.8150 ;
      RECT 3.2300 1.4200 3.3200 1.7250 ;
      RECT 3.2300 1.3300 3.3500 1.4200 ;
      RECT 3.2600 0.7200 3.3500 1.3300 ;
      RECT 2.9100 0.6300 3.3500 0.7200 ;
      RECT 2.2050 0.4300 2.3950 0.5100 ;
      RECT 2.9100 0.6000 3.0000 0.6300 ;
      RECT 2.3050 0.5200 3.0000 0.6000 ;
      RECT 2.2050 0.5100 3.0000 0.5200 ;
  END
END PREICG_X1B_A12TH

MACRO PREICG_X1P2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6650 ;
        RECT 0.8800 0.3200 0.9800 0.5700 ;
        RECT 1.9700 0.3200 2.0700 0.6300 ;
        RECT 3.0350 0.3200 3.1350 0.6550 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9500 1.5500 ;
        RECT 0.8500 1.5500 0.9500 1.6400 ;
        RECT 0.2500 0.8600 0.3500 1.4500 ;
        RECT 0.8500 1.6400 1.8250 1.7400 ;
        RECT 1.7250 1.3250 1.8250 1.6400 ;
        RECT 1.3350 0.9650 1.4250 1.6400 ;
        RECT 1.7250 1.2350 2.4900 1.3250 ;
        RECT 1.3350 0.8750 1.6000 0.9650 ;
        RECT 2.4000 1.1150 2.4900 1.2350 ;
        RECT 1.5100 0.6900 1.6000 0.8750 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5000 1.0500 0.9600 1.1500 ;
    END
    ANTENNAGATEAREA 0.0432 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5900 0.8500 1.0100 0.9500 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END E

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1650 1.4500 3.5500 1.5500 ;
        RECT 3.1650 1.5500 3.2650 1.9800 ;
        RECT 3.4500 0.7800 3.5500 1.4500 ;
        RECT 3.2950 0.6800 3.5500 0.7800 ;
        RECT 3.2950 0.4100 3.3950 0.6800 ;
    END
    ANTENNADIFFAREA 0.2071 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 2.9050 1.7750 3.0050 2.0800 ;
        RECT 2.2750 1.7700 2.3650 2.0800 ;
        RECT 3.4250 1.7550 3.5250 2.0800 ;
        RECT 1.9150 1.5150 2.0150 2.0800 ;
        RECT 1.9150 1.4150 2.1250 1.5150 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2350 1.4150 2.7600 1.5050 ;
      RECT 2.6700 0.9650 2.7600 1.4150 ;
      RECT 1.8700 0.8750 2.7600 0.9650 ;
      RECT 2.2350 1.5050 2.3250 1.6050 ;
      RECT 2.2350 0.4400 2.3250 0.8750 ;
      RECT 1.8700 0.7650 1.9600 0.8750 ;
      RECT 2.8500 1.2700 3.2850 1.3600 ;
      RECT 3.1950 0.9400 3.2850 1.2700 ;
      RECT 2.5550 1.5950 2.9400 1.6850 ;
      RECT 2.8500 1.3600 2.9400 1.5950 ;
      RECT 2.8500 0.7800 2.9400 1.2700 ;
      RECT 2.4950 0.6900 2.9400 0.7800 ;
      RECT 2.5550 1.6850 2.6450 1.9700 ;
      RECT 2.4950 0.4100 2.5850 0.6900 ;
      RECT 1.0550 1.4100 1.2450 1.5000 ;
      RECT 1.1550 0.7500 1.2450 1.4100 ;
      RECT 0.6200 0.6600 1.2450 0.7500 ;
      RECT 1.1550 0.4300 1.2450 0.6600 ;
      RECT 0.6200 0.4400 0.7100 0.6600 ;
      RECT 0.6600 1.8300 1.7700 1.9200 ;
      RECT 0.6600 1.7400 0.7500 1.8300 ;
      RECT 0.0700 1.6500 0.7500 1.7400 ;
      RECT 0.0700 1.7400 0.1700 1.8650 ;
      RECT 0.0700 0.6700 0.1600 1.6500 ;
      RECT 0.0700 0.4700 0.2050 0.6700 ;
      RECT 1.5150 1.0550 2.2800 1.1450 ;
      RECT 1.6900 0.5800 1.7800 1.0550 ;
      RECT 1.3850 0.4900 1.7800 0.5800 ;
      RECT 1.5150 1.1450 1.6050 1.5300 ;
  END
END PREICG_X1P2B_A12TH

MACRO PREICG_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3600 0.3200 0.4600 0.6050 ;
        RECT 0.8800 0.3200 0.9800 0.5200 ;
        RECT 1.9950 0.3200 2.0950 0.6200 ;
        RECT 3.1200 0.3200 3.2200 0.6050 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8300 0.3500 1.4500 ;
        RECT 0.2500 1.4500 0.9650 1.5500 ;
        RECT 0.8650 1.5500 0.9650 1.6400 ;
        RECT 0.8650 1.6400 1.8500 1.7400 ;
        RECT 1.7600 1.2850 1.8500 1.6400 ;
        RECT 1.3250 0.8700 1.4150 1.6400 ;
        RECT 1.7600 1.1950 2.5450 1.2850 ;
        RECT 1.3250 0.7800 1.6150 0.8700 ;
        RECT 2.4550 1.0700 2.5450 1.1950 ;
        RECT 1.5250 0.6900 1.6150 0.7800 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8400 1.0450 0.9500 ;
    END
    ANTENNAGATEAREA 0.0351 ;
  END E

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1550 1.4500 3.5500 1.5500 ;
        RECT 3.1550 1.5500 3.2550 1.9750 ;
        RECT 3.4500 0.8850 3.5500 1.4500 ;
        RECT 3.4100 0.4550 3.5500 0.8850 ;
    END
    ANTENNADIFFAREA 0.23495 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 2.8200 1.7750 3.0000 2.0800 ;
        RECT 2.2950 1.7500 2.3950 2.0800 ;
        RECT 3.4250 1.7500 3.5250 2.0800 ;
        RECT 2.0300 1.4750 2.1300 2.0800 ;
        RECT 1.9600 1.3750 2.1300 1.4750 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2600 1.3950 2.8300 1.4850 ;
      RECT 2.7400 0.9250 2.8300 1.3950 ;
      RECT 1.8900 0.8350 2.8300 0.9250 ;
      RECT 2.2600 1.4850 2.3500 1.5850 ;
      RECT 2.2600 0.4300 2.3600 0.8350 ;
      RECT 1.8900 0.7300 1.9800 0.8350 ;
      RECT 2.9400 1.1900 3.3600 1.2800 ;
      RECT 2.5600 1.5750 3.0300 1.6650 ;
      RECT 2.9400 1.2800 3.0300 1.5750 ;
      RECT 2.9400 0.7450 3.0300 1.1900 ;
      RECT 2.6250 0.6550 3.0300 0.7450 ;
      RECT 2.5600 1.6650 2.6500 1.9550 ;
      RECT 2.6250 0.4500 2.7150 0.6550 ;
      RECT 1.1350 0.7000 1.2250 1.5300 ;
      RECT 0.6250 0.6100 1.2250 0.7000 ;
      RECT 1.1350 0.4100 1.2250 0.6100 ;
      RECT 0.6250 0.4250 0.7150 0.6100 ;
      RECT 0.6850 1.8300 1.7600 1.9200 ;
      RECT 0.0450 1.7400 0.1700 1.8400 ;
      RECT 0.0450 0.6200 0.1450 1.6500 ;
      RECT 0.0450 0.4100 0.1700 0.6200 ;
      RECT 0.6850 1.7400 0.7750 1.8300 ;
      RECT 0.0450 1.6500 0.7750 1.7400 ;
      RECT 1.5050 1.0150 2.2550 1.1050 ;
      RECT 1.7100 0.5800 1.8000 1.0150 ;
      RECT 1.3350 0.4900 1.8000 0.5800 ;
      RECT 1.5050 1.1050 1.5950 1.5300 ;
  END
END PREICG_X1P4B_A12TH

MACRO PREICG_X1P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.6300 ;
        RECT 0.9250 0.3200 1.0250 0.5700 ;
        RECT 2.0100 0.3200 2.1100 0.5950 ;
        RECT 3.0550 0.3200 3.1550 0.5800 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8900 1.2500 2.6950 1.3500 ;
        RECT 1.8900 1.3500 1.9900 1.6400 ;
        RECT 2.5950 1.0500 2.6950 1.2500 ;
        RECT 0.7300 1.6400 1.9900 1.7400 ;
        RECT 0.7300 1.4950 0.8300 1.6400 ;
        RECT 1.2400 1.3250 1.3400 1.6400 ;
        RECT 0.2600 1.3950 0.8300 1.4950 ;
        RECT 1.2400 1.2250 1.6100 1.3250 ;
        RECT 0.2600 1.1000 0.3500 1.3950 ;
        RECT 1.5100 0.7000 1.6100 1.2250 ;
    END
    ANTENNAGATEAREA 0.1074 ;
  END CK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 0.8500 0.7050 0.9500 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.0500 0.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0372 ;
  END E

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3650 1.4500 3.7500 1.5500 ;
        RECT 3.3650 1.5500 3.4650 1.8800 ;
        RECT 3.6500 0.9500 3.7500 1.4500 ;
        RECT 3.3600 0.8500 3.7500 0.9500 ;
        RECT 3.3600 0.5100 3.4600 0.8500 ;
    END
    ANTENNADIFFAREA 0.3399 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.3350 1.7850 0.4350 2.0800 ;
        RECT 3.6250 1.7750 3.7250 2.0800 ;
        RECT 2.4250 1.7700 2.5250 2.0800 ;
        RECT 2.0800 1.4700 2.2500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6600 0.6600 1.2750 0.7500 ;
      RECT 1.1850 0.4100 1.2750 0.6600 ;
      RECT 0.9400 1.4450 1.1500 1.5450 ;
      RECT 1.0600 0.7500 1.1500 1.4450 ;
      RECT 0.6600 0.4300 0.7500 0.6600 ;
      RECT 0.5400 1.8300 1.7650 1.9200 ;
      RECT 0.0800 1.6750 0.1700 1.9650 ;
      RECT 0.0800 0.4350 0.1700 1.5850 ;
      RECT 0.5400 1.6750 0.6300 1.8300 ;
      RECT 0.0800 1.5850 0.6300 1.6750 ;
      RECT 1.7000 1.0500 2.3750 1.1400 ;
      RECT 1.4500 1.4400 1.7900 1.5300 ;
      RECT 1.7000 1.1400 1.7900 1.4400 ;
      RECT 1.7000 0.5500 1.7900 1.0500 ;
      RECT 1.3850 0.4600 1.7900 0.5500 ;
      RECT 2.3600 1.4400 2.9700 1.5300 ;
      RECT 2.8800 0.9600 2.9700 1.4400 ;
      RECT 1.8850 0.8700 2.9700 0.9600 ;
      RECT 2.2250 0.5200 2.3150 0.8700 ;
      RECT 2.2250 0.4300 2.4050 0.5200 ;
      RECT 1.8850 0.7500 1.9750 0.8700 ;
      RECT 3.1650 1.1750 3.5100 1.2650 ;
      RECT 2.6350 1.8050 3.2550 1.8950 ;
      RECT 3.1650 1.2650 3.2550 1.8050 ;
      RECT 3.1650 0.7800 3.2550 1.1750 ;
      RECT 2.5150 0.6900 3.2550 0.7800 ;
      RECT 2.5150 0.5050 2.6050 0.6900 ;
  END
END PREICG_X1P7B_A12TH

MACRO PREICG_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5300 ;
        RECT 0.5950 0.3200 0.6950 0.5750 ;
        RECT 2.0400 0.3200 2.1450 0.6600 ;
        RECT 3.1050 0.3200 3.2050 0.7100 ;
        RECT 3.6250 0.3200 3.7250 0.7100 ;
    END
  END VSS

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9650 0.1600 1.3650 ;
    END
    ANTENNAGATEAREA 0.0393 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9100 0.5500 1.3950 ;
    END
    ANTENNAGATEAREA 0.0507 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.3150 0.7500 1.8200 ;
        RECT 0.6500 1.8200 1.7500 1.9200 ;
        RECT 0.6500 1.2250 0.8750 1.3150 ;
        RECT 1.6500 1.4550 1.7500 1.8200 ;
        RECT 0.7750 0.8750 0.8750 1.2250 ;
        RECT 1.6500 1.3550 2.7900 1.4550 ;
        RECT 2.6850 1.2450 2.7900 1.3550 ;
    END
    ANTENNAGATEAREA 0.1173 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3650 1.2500 3.7500 1.3500 ;
        RECT 3.3650 1.3500 3.4650 1.7200 ;
        RECT 3.6500 0.9500 3.7500 1.2500 ;
        RECT 3.3650 0.8500 3.7500 0.9500 ;
        RECT 3.3650 0.5250 3.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.6050 2.0100 0.7050 2.0800 ;
        RECT 2.4700 1.9350 2.5700 2.0800 ;
        RECT 3.6250 1.7700 3.7250 2.0800 ;
        RECT 1.9850 1.5950 2.0850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2500 0.6800 1.1550 0.7700 ;
      RECT 1.0650 0.7700 1.1550 1.5250 ;
      RECT 0.0800 1.6800 0.1700 1.9800 ;
      RECT 0.0800 1.5900 0.3400 1.6800 ;
      RECT 0.2500 0.7700 0.3400 1.5900 ;
      RECT 0.3400 0.4100 0.4300 0.6800 ;
      RECT 1.2450 0.9950 1.8150 1.0850 ;
      RECT 0.9100 1.6400 1.3350 1.7300 ;
      RECT 1.2450 1.0850 1.3350 1.6400 ;
      RECT 1.2450 0.5900 1.3350 0.9950 ;
      RECT 0.9650 0.5250 1.3350 0.5900 ;
      RECT 0.8250 0.5000 1.3350 0.5250 ;
      RECT 0.8250 0.4350 1.0550 0.5000 ;
      RECT 1.8200 0.7900 2.3050 0.8800 ;
      RECT 1.4250 1.1750 2.0150 1.2650 ;
      RECT 1.9250 0.8800 2.0150 1.1750 ;
      RECT 1.8200 0.6800 1.9100 0.7900 ;
      RECT 1.4250 0.5900 1.9100 0.6800 ;
      RECT 1.4250 1.2650 1.5150 1.5700 ;
      RECT 1.4250 0.4700 1.5150 0.5900 ;
      RECT 2.2300 1.6050 3.0600 1.6950 ;
      RECT 2.9700 1.1200 3.0600 1.6050 ;
      RECT 2.1050 1.0300 3.0600 1.1200 ;
      RECT 2.1050 1.1200 2.1950 1.2400 ;
      RECT 2.4150 0.6000 2.5050 1.0300 ;
      RECT 2.2550 0.5100 2.5050 0.6000 ;
      RECT 3.1600 1.0450 3.5400 1.1350 ;
      RECT 2.6750 1.8100 3.2500 1.9000 ;
      RECT 3.1600 1.1350 3.2500 1.8100 ;
      RECT 3.1600 0.9400 3.2500 1.0450 ;
      RECT 2.6150 0.8500 3.2500 0.9400 ;
      RECT 2.6150 0.4400 2.7050 0.8500 ;
  END
END PREICG_X2B_A12TH

MACRO PREICG_X2P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7200 ;
        RECT 2.4150 0.3200 2.6350 0.3700 ;
        RECT 3.2450 0.3200 3.3450 0.9200 ;
        RECT 3.7650 0.3200 3.8650 0.7150 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.0900 1.7250 0.1900 2.0800 ;
        RECT 2.9950 1.6700 3.0950 2.0800 ;
        RECT 3.2450 1.6250 3.3450 2.0800 ;
        RECT 3.7650 1.6250 3.8650 2.0800 ;
        RECT 2.4750 1.3350 2.5750 2.0800 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4950 ;
    END
    ANTENNAGATEAREA 0.0555 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1050 0.5500 1.5750 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.5700 1.3500 0.9900 ;
        RECT 0.8200 0.4800 2.9100 0.5700 ;
        RECT 0.8200 0.5700 0.9100 1.4700 ;
        RECT 2.1750 0.5700 2.3450 0.5800 ;
        RECT 2.8100 0.5700 2.9100 1.2650 ;
    END
    ANTENNAGATEAREA 0.1344 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.9500 4.1500 1.2500 ;
        RECT 3.5050 1.2500 4.1500 1.3500 ;
        RECT 3.5050 0.8500 4.1500 0.9500 ;
        RECT 3.5050 1.3500 3.6050 1.6900 ;
        RECT 4.0300 1.3500 4.1500 1.6900 ;
        RECT 3.5050 0.5050 3.6050 0.8500 ;
        RECT 4.0250 0.5050 4.1500 0.8500 ;
    END
    ANTENNADIFFAREA 0.4086 ;
  END ECK
  OBS
    LAYER M1 ;
      RECT 0.6400 0.9000 0.7300 1.7450 ;
      RECT 0.0950 0.8100 0.7300 0.9000 ;
      RECT 0.6400 0.6200 0.7300 0.8100 ;
      RECT 0.0950 0.6200 0.1850 0.8100 ;
      RECT 1.0200 1.1250 1.7450 1.2150 ;
      RECT 1.6550 1.0100 1.7450 1.1250 ;
      RECT 0.8600 1.5800 1.1100 1.6700 ;
      RECT 1.0200 1.2150 1.1100 1.5800 ;
      RECT 1.0200 0.6900 1.1100 1.1250 ;
      RECT 1.0300 1.8450 1.3200 1.9350 ;
      RECT 1.2300 1.8400 1.3200 1.8450 ;
      RECT 1.2300 1.7500 2.2300 1.8400 ;
      RECT 2.1400 0.9400 2.2300 1.7500 ;
      RECT 2.0600 0.8500 2.2300 0.9400 ;
      RECT 1.8500 0.6700 2.6450 0.7600 ;
      RECT 2.5550 0.7600 2.6450 1.2150 ;
      RECT 1.8250 1.3950 1.9950 1.6550 ;
      RECT 1.2600 1.3050 1.9950 1.3950 ;
      RECT 1.8500 0.7600 1.9400 1.3050 ;
      RECT 3.0000 1.0550 3.8950 1.1450 ;
      RECT 2.6850 1.3950 3.0900 1.4850 ;
      RECT 3.0000 1.1450 3.0900 1.3950 ;
      RECT 3.0000 0.5600 3.0900 1.0550 ;
  END
END PREICG_X2P5B_A12TH

MACRO PREICG_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.6100 ;
        RECT 2.3900 0.3200 2.5600 0.3900 ;
        RECT 3.4200 0.3200 3.5200 0.7100 ;
        RECT 3.9650 0.3200 4.0650 0.7350 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.9100 0.3550 1.3050 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0450 0.5500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0471 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0500 3.1450 1.1500 ;
        RECT 2.6500 0.5800 2.7500 1.0500 ;
        RECT 0.8200 0.4800 2.7500 0.5800 ;
        RECT 0.8200 0.5800 0.9200 1.4700 ;
    END
    ANTENNAGATEAREA 0.1518 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9550 4.3500 1.2500 ;
        RECT 3.7050 1.2500 4.3500 1.3500 ;
        RECT 3.7050 0.8550 4.3500 0.9550 ;
        RECT 3.7050 1.3500 3.8050 1.7200 ;
        RECT 4.2300 1.3500 4.3500 1.7200 ;
        RECT 3.7050 0.5350 3.8050 0.8550 ;
        RECT 4.2300 0.5350 4.3500 0.8550 ;
    END
    ANTENNADIFFAREA 0.4914 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 3.4450 1.7700 3.5450 2.0800 ;
        RECT 3.9650 1.7700 4.0650 2.0800 ;
        RECT 2.7800 1.6800 2.8800 2.0800 ;
        RECT 1.4800 1.6650 1.5800 2.0800 ;
        RECT 0.0900 1.6600 0.1900 2.0800 ;
        RECT 2.2700 1.5350 2.3700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6400 0.8200 0.7300 1.9000 ;
      RECT 0.0950 0.7300 0.7300 0.8200 ;
      RECT 0.6400 0.6200 0.7300 0.7300 ;
      RECT 0.0950 0.6200 0.1850 0.7300 ;
      RECT 1.0550 1.0750 1.7900 1.1650 ;
      RECT 0.8400 1.5800 1.1450 1.6700 ;
      RECT 1.0550 1.1650 1.1450 1.5800 ;
      RECT 1.0550 0.8650 1.1450 1.0750 ;
      RECT 1.0200 0.6950 1.1450 0.8650 ;
      RECT 2.0850 0.8500 2.2750 0.9400 ;
      RECT 1.0300 1.8450 1.3450 1.9350 ;
      RECT 1.2550 1.5750 1.3450 1.8450 ;
      RECT 1.2550 1.4850 2.1750 1.5750 ;
      RECT 2.0150 1.5750 2.1050 1.7450 ;
      RECT 2.0850 0.9400 2.1750 1.4850 ;
      RECT 2.4500 1.3000 3.3950 1.3900 ;
      RECT 1.2650 1.3050 1.9700 1.3950 ;
      RECT 1.8800 0.7600 1.9700 1.3050 ;
      RECT 1.8800 0.6700 2.5400 0.7600 ;
      RECT 2.4500 0.7600 2.5400 1.0450 ;
      RECT 2.4500 1.0450 2.5500 1.3000 ;
      RECT 3.5000 1.0500 4.1000 1.1500 ;
      RECT 3.0700 1.5900 3.1700 1.7800 ;
      RECT 2.9400 0.5150 3.0300 0.8150 ;
      RECT 2.5200 1.5000 3.5900 1.5900 ;
      RECT 3.5000 1.1500 3.5900 1.5000 ;
      RECT 3.5000 0.9050 3.5900 1.0500 ;
      RECT 2.9400 0.8150 3.5900 0.9050 ;
      RECT 2.5200 1.5900 2.6200 1.9800 ;
  END
END PREICG_X3B_A12TH

MACRO PREICG_X3P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.6100 ;
        RECT 2.3900 0.3200 2.5600 0.3900 ;
        RECT 3.3850 0.3200 3.4850 0.7200 ;
        RECT 3.9050 0.3200 4.0050 0.7500 ;
        RECT 4.4250 0.3200 4.5250 0.7500 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9550 4.3500 1.2500 ;
        RECT 3.6450 1.2500 4.3500 1.3500 ;
        RECT 3.6450 0.8550 4.3500 0.9550 ;
        RECT 3.6450 1.3500 3.7450 1.7200 ;
        RECT 4.1650 1.3500 4.2650 1.7200 ;
        RECT 3.6450 0.5350 3.7450 0.8550 ;
        RECT 4.1650 0.5350 4.2650 0.8550 ;
    END
    ANTENNADIFFAREA 0.478 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0500 3.1350 1.1500 ;
        RECT 2.6500 0.5800 2.7500 1.0500 ;
        RECT 0.8200 0.4800 2.7500 0.5800 ;
        RECT 0.8200 0.5800 0.9200 1.4700 ;
    END
    ANTENNAGATEAREA 0.1689 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 3.3750 1.9050 3.4950 2.0800 ;
        RECT 0.0900 1.7100 0.1900 2.0800 ;
        RECT 2.7700 1.7000 2.8700 2.0800 ;
        RECT 4.4250 1.6800 4.5250 2.0800 ;
        RECT 1.4800 1.6650 1.5800 2.0800 ;
        RECT 3.9050 1.6650 4.0050 2.0800 ;
        RECT 2.2250 1.6500 2.3950 2.0800 ;
    END
  END VDD

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0450 0.5500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0507 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.9100 0.3550 1.3050 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 3.2350 1.3900 3.3250 1.4300 ;
      RECT 2.4400 1.3000 3.3250 1.3900 ;
      RECT 3.2350 1.2600 3.3250 1.3000 ;
      RECT 2.4400 1.0500 2.5500 1.3000 ;
      RECT 2.4400 0.7600 2.5300 1.0500 ;
      RECT 1.8800 0.6700 2.5300 0.7600 ;
      RECT 1.8800 0.7600 1.9700 1.3050 ;
      RECT 1.2650 1.3050 1.9700 1.3950 ;
      RECT 3.4450 1.0500 4.0400 1.1500 ;
      RECT 3.0500 1.6100 3.1500 1.7350 ;
      RECT 2.9250 0.4900 3.0250 0.8100 ;
      RECT 2.5100 1.5200 3.5350 1.6100 ;
      RECT 3.4450 1.1500 3.5350 1.5200 ;
      RECT 3.4450 0.9000 3.5350 1.0500 ;
      RECT 2.9250 0.8100 3.5350 0.9000 ;
      RECT 2.5100 1.6100 2.6100 1.9850 ;
      RECT 0.6400 0.8200 0.7300 1.9000 ;
      RECT 0.0550 0.7300 0.7300 0.8200 ;
      RECT 0.6400 0.4600 0.7300 0.7300 ;
      RECT 0.0550 0.4950 0.2250 0.7300 ;
      RECT 1.0550 1.0750 1.7900 1.1650 ;
      RECT 0.8400 1.5800 1.1450 1.6700 ;
      RECT 1.0550 1.1650 1.1450 1.5800 ;
      RECT 1.0550 0.8650 1.1450 1.0750 ;
      RECT 1.0200 0.6950 1.1450 0.8650 ;
      RECT 2.0850 0.8500 2.2550 0.9400 ;
      RECT 1.0100 1.8450 1.3500 1.9350 ;
      RECT 1.2600 1.5750 1.3500 1.8450 ;
      RECT 1.2600 1.4850 2.1750 1.5750 ;
      RECT 2.0050 1.5750 2.0950 1.7800 ;
      RECT 2.0850 0.9400 2.1750 1.4850 ;
  END
END PREICG_X3P5B_A12TH

MACRO PREICG_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6400 ;
        RECT 2.3900 0.3200 2.5600 0.3900 ;
        RECT 3.3850 0.3200 3.4850 0.6900 ;
        RECT 3.9050 0.3200 4.0050 0.7050 ;
        RECT 4.4250 0.3200 4.5250 0.7000 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9550 4.3500 1.2500 ;
        RECT 3.6450 1.2500 4.3500 1.3500 ;
        RECT 3.6450 0.8550 4.3500 0.9550 ;
        RECT 3.6450 1.3500 3.7450 1.7200 ;
        RECT 4.1650 1.3500 4.2650 1.7200 ;
        RECT 3.6450 0.5350 3.7450 0.8550 ;
        RECT 4.1650 0.5350 4.2650 0.8550 ;
    END
    ANTENNADIFFAREA 0.546 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0500 3.1350 1.1500 ;
        RECT 2.6500 0.5800 2.7500 1.0500 ;
        RECT 0.8200 0.4800 2.7500 0.5800 ;
        RECT 0.8200 0.5800 0.9200 1.4700 ;
    END
    ANTENNAGATEAREA 0.1857 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0450 0.5500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.9100 0.3550 1.3050 ;
    END
    ANTENNAGATEAREA 0.0702 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 3.3850 1.8600 3.4850 2.0800 ;
        RECT 3.9050 1.7750 4.0050 2.0800 ;
        RECT 4.4250 1.7750 4.5250 2.0800 ;
        RECT 0.0900 1.7400 0.1900 2.0800 ;
        RECT 2.7700 1.7000 2.8700 2.0800 ;
        RECT 1.4800 1.6650 1.5800 2.0800 ;
        RECT 2.2250 1.6500 2.3950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.4400 1.3400 3.3250 1.4300 ;
      RECT 3.2350 1.2600 3.3250 1.3400 ;
      RECT 1.2650 1.3050 1.9700 1.3950 ;
      RECT 1.8800 0.7600 1.9700 1.3050 ;
      RECT 1.8800 0.6700 2.5300 0.7600 ;
      RECT 2.4400 0.7600 2.5300 1.0500 ;
      RECT 2.4400 1.0500 2.5500 1.3400 ;
      RECT 3.4450 1.0500 4.0400 1.1500 ;
      RECT 3.0500 1.6100 3.1500 1.7350 ;
      RECT 2.9250 0.4700 3.0250 0.8100 ;
      RECT 2.5100 1.5200 3.5350 1.6100 ;
      RECT 3.4450 1.1500 3.5350 1.5200 ;
      RECT 3.4450 0.9000 3.5350 1.0500 ;
      RECT 2.9250 0.8100 3.5350 0.9000 ;
      RECT 2.5100 1.6100 2.6100 1.9850 ;
      RECT 0.6400 0.8200 0.7300 1.9000 ;
      RECT 0.0950 0.7300 0.7300 0.8200 ;
      RECT 0.6400 0.4600 0.7300 0.7300 ;
      RECT 0.0950 0.4300 0.1850 0.7300 ;
      RECT 1.0550 1.0750 1.7900 1.1650 ;
      RECT 0.8400 1.5800 1.1450 1.6700 ;
      RECT 1.0550 1.1650 1.1450 1.5800 ;
      RECT 1.0550 0.8650 1.1450 1.0750 ;
      RECT 1.0200 0.6950 1.1450 0.8650 ;
      RECT 2.0850 0.8500 2.2550 0.9400 ;
      RECT 1.0100 1.8450 1.3550 1.9350 ;
      RECT 1.2650 1.5750 1.3550 1.8450 ;
      RECT 1.2650 1.4850 2.1750 1.5750 ;
      RECT 2.0050 1.5750 2.0950 1.7800 ;
      RECT 2.0850 0.9400 2.1750 1.4850 ;
  END
END PREICG_X4B_A12TH

MACRO PREICG_X5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.7150 ;
        RECT 3.4150 0.3200 3.5150 0.6300 ;
        RECT 4.0450 0.3200 4.1450 0.6950 ;
        RECT 4.5650 0.3200 4.6650 0.6950 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 3.5250 1.7700 3.6250 2.0800 ;
        RECT 4.0450 1.7650 4.1450 2.0800 ;
        RECT 4.5650 1.7650 4.6650 2.0800 ;
        RECT 1.4600 1.6650 1.5600 2.0800 ;
        RECT 2.8550 1.5350 2.9550 2.0800 ;
        RECT 2.3050 1.3500 2.4050 2.0800 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.1000 0.3500 1.3050 ;
        RECT 0.0950 1.0000 0.3500 1.1000 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.5050 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.5800 2.7500 0.9650 ;
        RECT 2.6500 0.9650 3.1350 1.0650 ;
        RECT 0.8200 0.4800 2.7500 0.5800 ;
        RECT 0.8200 0.5800 0.9200 1.4700 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8300 0.9500 4.9500 1.2500 ;
        RECT 3.7850 1.2500 4.9500 1.3500 ;
        RECT 3.7850 0.8500 4.9500 0.9500 ;
        RECT 3.7850 1.3500 3.8850 1.7000 ;
        RECT 4.3050 1.3500 4.4050 1.7000 ;
        RECT 4.8300 1.3500 4.9500 1.7000 ;
        RECT 3.7850 0.5400 3.8850 0.8500 ;
        RECT 4.3050 0.5400 4.4050 0.8500 ;
        RECT 4.8300 0.5400 4.9500 0.8500 ;
    END
    ANTENNADIFFAREA 0.8344 ;
  END ECK
  OBS
    LAYER M1 ;
      RECT 0.6400 0.9000 0.7300 1.9300 ;
      RECT 0.0950 0.8100 0.7300 0.9000 ;
      RECT 0.6400 0.4400 0.7300 0.8100 ;
      RECT 0.0950 0.4400 0.1850 0.8100 ;
      RECT 1.0550 1.0750 1.7350 1.1650 ;
      RECT 0.8400 1.5800 1.1450 1.6700 ;
      RECT 1.0550 1.1650 1.1450 1.5800 ;
      RECT 1.0550 0.8600 1.1450 1.0750 ;
      RECT 1.0100 0.6900 1.1450 0.8600 ;
      RECT 1.2550 1.4850 2.1400 1.5750 ;
      RECT 2.0500 0.9400 2.1400 1.4850 ;
      RECT 2.0500 0.8500 2.2350 0.9400 ;
      RECT 1.0000 1.8450 1.3450 1.9350 ;
      RECT 1.2550 1.5750 1.3450 1.8450 ;
      RECT 2.4550 1.1550 3.4000 1.2450 ;
      RECT 3.3100 0.9850 3.4000 1.1550 ;
      RECT 1.7350 0.6700 2.5450 0.7600 ;
      RECT 2.4550 0.7600 2.5450 1.0400 ;
      RECT 2.4550 1.0400 2.5500 1.1550 ;
      RECT 1.2600 1.3050 1.9150 1.3950 ;
      RECT 1.8250 0.7600 1.9150 1.3050 ;
      RECT 3.5100 1.0500 4.5000 1.1500 ;
      RECT 2.8600 0.4500 2.9500 0.7850 ;
      RECT 2.6000 1.4250 2.6900 1.7500 ;
      RECT 2.6000 1.3350 3.6000 1.4250 ;
      RECT 3.5100 1.1500 3.6000 1.3350 ;
      RECT 3.5100 0.8750 3.6000 1.0500 ;
      RECT 2.8600 0.7850 3.6000 0.8750 ;
  END
END PREICG_X5B_A12TH

MACRO PREICG_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.4850 0.3200 0.5850 0.7100 ;
        RECT 3.6200 0.3200 3.7900 0.6300 ;
        RECT 4.1850 0.3200 4.2850 0.7250 ;
        RECT 4.7050 0.3200 4.8050 0.7250 ;
        RECT 5.2250 0.3200 5.3250 0.7200 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0850 0.3550 1.4850 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END SE

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6550 1.2550 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9950 1.0350 3.4450 1.1500 ;
        RECT 2.9950 0.5800 3.0950 1.0350 ;
        RECT 0.9350 0.4800 3.0950 0.5800 ;
        RECT 0.9350 0.5800 1.0350 1.3400 ;
        RECT 0.9350 1.3400 1.1500 1.4300 ;
    END
    ANTENNAGATEAREA 0.2496 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.9500 5.1500 1.2500 ;
        RECT 3.9250 1.2500 5.1500 1.3500 ;
        RECT 3.9250 0.8500 5.1500 0.9500 ;
        RECT 3.9250 1.3500 4.0250 1.7200 ;
        RECT 4.4450 1.3500 4.5450 1.7200 ;
        RECT 4.9650 1.3500 5.0650 1.7200 ;
        RECT 3.9250 0.5200 4.0250 0.8500 ;
        RECT 4.4450 0.5200 4.5450 0.8500 ;
        RECT 4.9650 0.5200 5.0650 0.8500 ;
    END
    ANTENNADIFFAREA 0.894 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 0.3000 1.9300 0.4700 2.0800 ;
        RECT 3.6650 1.8100 3.7650 2.0800 ;
        RECT 3.0550 1.8000 3.1550 2.0800 ;
        RECT 4.1850 1.7700 4.2850 2.0800 ;
        RECT 4.7050 1.7700 4.8050 2.0800 ;
        RECT 5.2250 1.7700 5.3250 2.0800 ;
        RECT 2.1750 1.6800 2.3450 2.0800 ;
        RECT 1.6850 1.6650 1.7850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.7500 0.7500 1.8400 ;
      RECT 0.0750 1.8400 0.1750 1.9600 ;
      RECT 0.8650 1.6300 0.9550 1.9650 ;
      RECT 0.7550 1.5400 0.9550 1.6300 ;
      RECT 0.7550 0.8900 0.8450 1.5400 ;
      RECT 0.2300 0.8000 0.8450 0.8900 ;
      RECT 0.7550 0.4400 0.8450 0.8000 ;
      RECT 0.2300 0.4600 0.3200 0.8000 ;
      RECT 1.2800 1.0750 2.1700 1.1650 ;
      RECT 1.0850 1.5800 1.3700 1.6700 ;
      RECT 1.2800 1.1650 1.3700 1.5800 ;
      RECT 1.2800 0.9050 1.3700 1.0750 ;
      RECT 1.1250 0.8150 1.3700 0.9050 ;
      RECT 1.1250 0.6950 1.2150 0.8150 ;
      RECT 1.4850 1.4850 2.6400 1.5750 ;
      RECT 2.5500 0.9400 2.6400 1.4850 ;
      RECT 2.4950 0.8500 2.6650 0.9400 ;
      RECT 1.2400 1.8450 1.5750 1.9350 ;
      RECT 1.4850 1.5750 1.5750 1.8450 ;
      RECT 2.7950 1.2800 3.6350 1.3700 ;
      RECT 3.5450 1.0750 3.6350 1.2800 ;
      RECT 1.4850 1.3050 2.3500 1.3950 ;
      RECT 2.2600 0.7600 2.3500 1.3050 ;
      RECT 1.8350 0.6700 2.8850 0.7600 ;
      RECT 2.7950 0.7600 2.8850 1.2800 ;
      RECT 3.7450 1.0550 4.7150 1.1450 ;
      RECT 2.7950 1.5650 2.8950 1.9250 ;
      RECT 3.1850 0.4700 3.2850 0.8100 ;
      RECT 2.7950 1.4750 3.8350 1.5650 ;
      RECT 3.7450 1.1450 3.8350 1.4750 ;
      RECT 3.7450 0.9000 3.8350 1.0550 ;
      RECT 3.1850 0.8100 3.8350 0.9000 ;
  END
END PREICG_X6B_A12TH

MACRO PREICG_X7P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.5400 ;
        RECT 3.5700 0.3200 3.6700 0.6200 ;
        RECT 4.3700 0.3200 4.4700 0.7250 ;
        RECT 4.8900 0.3200 4.9900 0.6400 ;
        RECT 5.4100 0.3200 5.5100 0.6400 ;
        RECT 5.9300 0.3200 6.0300 0.6400 ;
    END
  END VSS

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9950 0.5300 1.1900 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4050 0.3300 1.5900 ;
    END
    ANTENNAGATEAREA 0.1044 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8750 1.0500 4.0900 1.1500 ;
        RECT 2.8750 0.5800 2.9750 1.0500 ;
        RECT 0.8000 0.4800 2.9750 0.5800 ;
        RECT 0.8000 0.5800 0.9000 1.0050 ;
        RECT 1.0450 0.4650 1.2150 0.4800 ;
        RECT 0.8000 1.0050 1.1550 1.1050 ;
        RECT 1.0500 1.1050 1.1550 1.4550 ;
    END
    ANTENNAGATEAREA 0.3135 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8400 0.8650 5.9600 1.2500 ;
        RECT 4.3600 1.2500 6.0300 1.3700 ;
        RECT 4.6200 0.7450 5.9600 0.8650 ;
        RECT 4.3600 1.3700 4.4800 1.7800 ;
        RECT 4.8900 1.3700 4.9900 1.6800 ;
        RECT 5.4100 1.3700 5.5100 1.6800 ;
        RECT 5.9300 1.3700 6.0300 1.7800 ;
        RECT 4.6200 0.4300 4.7400 0.7450 ;
        RECT 5.1500 0.4300 5.2500 0.7450 ;
        RECT 5.6700 0.4300 5.7700 0.7450 ;
    END
    ANTENNADIFFAREA 1.1423 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.8500 1.7700 2.9500 2.0800 ;
        RECT 3.3700 1.7700 3.4700 2.0800 ;
        RECT 4.0700 1.7700 4.1700 2.0800 ;
        RECT 4.6300 1.7200 4.7300 2.0800 ;
        RECT 5.1500 1.7200 5.2500 2.0800 ;
        RECT 5.6700 1.7200 5.7700 2.0800 ;
        RECT 2.2650 1.7000 2.3650 2.0800 ;
        RECT 1.7250 1.6650 1.8250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.8300 0.7450 1.9200 ;
      RECT 0.8750 1.7100 0.9750 1.9900 ;
      RECT 0.6200 1.6200 0.9750 1.7100 ;
      RECT 0.6200 0.7400 0.7100 1.6200 ;
      RECT 0.0550 0.6500 0.7100 0.7400 ;
      RECT 0.6200 0.5300 0.7100 0.6500 ;
      RECT 0.0550 0.4500 0.2250 0.6500 ;
      RECT 1.2650 1.0750 2.0750 1.1650 ;
      RECT 1.1000 1.5800 1.3550 1.6700 ;
      RECT 1.2650 1.1650 1.3550 1.5800 ;
      RECT 1.2650 0.8850 1.3550 1.0750 ;
      RECT 1.0100 0.7950 1.3550 0.8850 ;
      RECT 1.0100 0.6700 1.1000 0.7950 ;
      RECT 1.4800 1.4850 2.7200 1.5750 ;
      RECT 2.4750 0.9400 2.5650 1.4850 ;
      RECT 2.3950 0.8500 2.5650 0.9400 ;
      RECT 1.2700 1.8250 1.5700 1.9150 ;
      RECT 1.4800 1.5750 1.5700 1.8250 ;
      RECT 2.6750 1.2600 3.7000 1.3500 ;
      RECT 1.5050 1.3050 2.2850 1.3950 ;
      RECT 2.1950 0.7600 2.2850 1.3050 ;
      RECT 1.7350 0.6700 2.7650 0.7600 ;
      RECT 2.6750 0.7600 2.7650 1.2600 ;
      RECT 4.1800 0.9750 5.6000 1.0750 ;
      RECT 3.1100 1.5900 3.2100 1.9800 ;
      RECT 3.1150 0.4500 3.2050 0.8100 ;
      RECT 3.8100 1.5900 3.9100 1.9800 ;
      RECT 3.1100 1.5000 4.2700 1.5900 ;
      RECT 4.1800 1.0750 4.2700 1.5000 ;
      RECT 4.1800 0.9000 4.2700 0.9750 ;
      RECT 3.1150 0.8100 4.2700 0.9000 ;
      RECT 4.0300 0.4450 4.1300 0.8100 ;
  END
END PREICG_X7P5B_A12TH

MACRO PREICG_X9B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.5950 0.3200 0.6950 0.6200 ;
        RECT 3.6450 0.3200 3.7450 0.7050 ;
        RECT 4.5950 0.3200 4.6950 0.7050 ;
        RECT 5.1900 0.3200 5.2900 0.6900 ;
        RECT 5.7100 0.3200 5.8100 0.6900 ;
        RECT 6.2300 0.3200 6.3300 0.6950 ;
        RECT 6.7500 0.3200 6.8500 0.6950 ;
    END
  END VSS

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9100 0.7700 1.3050 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0000 0.5050 1.1000 ;
        RECT 0.2500 1.1000 0.3500 1.3050 ;
    END
    ANTENNAGATEAREA 0.1182 ;
  END SE

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9500 1.0500 4.3650 1.1500 ;
        RECT 2.9500 0.5800 3.0500 1.0500 ;
        RECT 1.0550 0.4800 3.0500 0.5800 ;
        RECT 1.0550 0.5800 1.1550 1.4850 ;
    END
    ANTENNAGATEAREA 0.3666 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 4.6700 1.7700 4.7700 2.0800 ;
        RECT 5.1900 1.7700 5.2900 2.0800 ;
        RECT 5.7100 1.7700 5.8100 2.0800 ;
        RECT 6.2300 1.7700 6.3300 2.0800 ;
        RECT 6.7500 1.7700 6.8500 2.0800 ;
        RECT 0.3000 1.6750 0.4700 2.0800 ;
        RECT 1.6900 1.6700 1.8600 2.0800 ;
        RECT 3.1500 1.6450 3.2500 2.0800 ;
        RECT 3.8450 1.6450 3.9450 2.0800 ;
        RECT 4.3650 1.6450 4.4650 2.0800 ;
        RECT 2.6000 1.5200 2.6900 2.0800 ;
    END
  END VDD

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9300 1.2350 7.1100 1.3650 ;
        RECT 4.9300 1.3650 5.0300 1.7200 ;
        RECT 5.4500 1.3650 5.5500 1.7200 ;
        RECT 5.9700 1.3650 6.0700 1.7200 ;
        RECT 6.4900 1.3650 6.5900 1.7200 ;
        RECT 7.0100 1.3650 7.1100 1.7200 ;
        RECT 6.9800 0.9650 7.1100 1.2350 ;
        RECT 4.9300 0.8350 7.1100 0.9650 ;
        RECT 4.9300 0.5050 5.0300 0.8350 ;
        RECT 5.4500 0.5050 5.5500 0.8350 ;
        RECT 5.9700 0.5050 6.0700 0.8350 ;
        RECT 6.4900 0.5050 6.5900 0.8350 ;
        RECT 7.0100 0.4950 7.1100 0.8350 ;
    END
    ANTENNADIFFAREA 1.4304 ;
  END ECK
  OBS
    LAYER M1 ;
      RECT 0.0750 1.4800 0.7100 1.5800 ;
      RECT 0.6100 1.5800 0.7100 1.9100 ;
      RECT 0.0750 1.5800 0.1750 1.9100 ;
      RECT 0.8750 0.8000 0.9650 1.9550 ;
      RECT 0.3400 0.7100 0.9650 0.8000 ;
      RECT 0.8750 0.4300 0.9650 0.7100 ;
      RECT 0.3400 0.4100 0.4300 0.7100 ;
      RECT 1.2450 1.0800 1.9750 1.1700 ;
      RECT 1.8850 0.9800 1.9750 1.0800 ;
      RECT 1.0800 1.5950 1.3350 1.6850 ;
      RECT 1.2450 1.1700 1.3350 1.5950 ;
      RECT 1.2450 0.7050 1.3350 1.0800 ;
      RECT 1.4400 1.4900 2.4250 1.5800 ;
      RECT 2.3350 0.9400 2.4250 1.4900 ;
      RECT 2.2950 0.8500 2.4650 0.9400 ;
      RECT 1.2600 1.8450 1.5300 1.9350 ;
      RECT 1.4400 1.5800 1.5300 1.8450 ;
      RECT 2.7500 1.2400 4.5950 1.3300 ;
      RECT 1.5000 1.3100 2.1850 1.4000 ;
      RECT 2.0950 0.7600 2.1850 1.3100 ;
      RECT 2.0250 0.6700 2.8400 0.7600 ;
      RECT 2.7500 0.7600 2.8400 1.2400 ;
      RECT 4.7000 1.0550 6.7000 1.1450 ;
      RECT 2.8900 1.5300 2.9900 1.8800 ;
      RECT 3.4100 1.5300 3.5100 1.8800 ;
      RECT 3.1500 0.4700 3.2500 0.8100 ;
      RECT 4.1050 1.5300 4.2050 1.8800 ;
      RECT 4.1050 0.4700 4.2050 0.8100 ;
      RECT 2.8900 1.4400 4.7900 1.5300 ;
      RECT 4.7000 1.1450 4.7900 1.4400 ;
      RECT 4.7000 0.9000 4.7900 1.0550 ;
      RECT 3.1500 0.8100 4.7900 0.9000 ;
  END
END PREICG_X9B_A12TH

MACRO RF1R1WS_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.4000 0.3200 0.5200 0.3900 ;
        RECT 1.6600 0.3200 1.7700 0.6850 ;
        RECT 1.9600 0.3200 2.1300 0.5400 ;
        RECT 3.0200 0.3200 3.1300 0.8800 ;
    END
  END VSS

  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9500 1.2100 3.1500 1.4250 ;
        RECT 2.9500 1.0300 3.0400 1.2100 ;
    END
    ANTENNAGATEAREA 0.0777 ;
  END RWL

  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.6200 0.9900 ;
        RECT 0.5300 0.9900 0.6200 1.3250 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END WBL

  PIN WWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.1900 0.3600 1.3900 ;
        RECT 0.2700 1.3900 0.3600 1.8000 ;
        RECT 0.2700 1.8000 1.2750 1.8900 ;
        RECT 1.1750 1.8900 1.2750 1.9800 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END WWL

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.4050 2.0400 0.5750 2.0800 ;
        RECT 1.9900 1.8100 2.1000 2.0800 ;
        RECT 3.0200 1.7900 3.1300 2.0800 ;
        RECT 1.5600 1.7600 1.6700 2.0800 ;
    END
  END VDD

  PIN RBL
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8900 2.5500 1.5850 ;
        RECT 2.4500 1.5850 2.6100 1.9550 ;
        RECT 2.4500 0.5200 2.6100 0.8900 ;
    END
    ANTENNADIFFAREA 0.2288 ;
  END RBL
  OBS
    LAYER M1 ;
      RECT 2.7700 1.4950 2.8600 1.9200 ;
      RECT 2.6950 1.3250 2.8600 1.4950 ;
      RECT 2.7700 0.7050 2.8600 1.3250 ;
      RECT 0.7200 0.6600 0.8100 1.6900 ;
      RECT 0.0550 0.4800 1.4150 0.5700 ;
      RECT 0.9200 0.5700 1.0100 1.4600 ;
      RECT 1.3250 0.5700 1.4150 1.0550 ;
      RECT 0.0550 1.5200 0.1750 1.8900 ;
      RECT 0.0550 0.7100 0.1450 1.5200 ;
      RECT 0.0550 0.5700 0.1950 0.7100 ;
      RECT 1.4400 1.3050 1.8300 1.3950 ;
      RECT 1.4400 1.2100 1.5400 1.3050 ;
      RECT 1.7400 0.9050 1.8300 1.3050 ;
      RECT 1.6350 0.8050 1.8300 0.9050 ;
      RECT 0.9400 1.5700 2.0650 1.6600 ;
      RECT 1.9750 1.0050 2.0650 1.5700 ;
      RECT 1.1200 0.6600 1.2100 1.5700 ;
      RECT 2.2600 0.5000 2.3500 1.9000 ;
  END
END RF1R1WS_X1M_A12TH

MACRO RF1R1WS_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 1.6300 0.3200 1.8000 0.4800 ;
        RECT 1.9400 0.3200 2.1100 0.5000 ;
        RECT 3.0800 0.3200 3.2900 0.3850 ;
    END
  END VSS

  PIN WWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.5900 2.7500 1.0950 ;
        RECT 2.6500 0.4900 3.3400 0.5900 ;
        RECT 3.2450 0.5900 3.3400 1.0650 ;
    END
    ANTENNAGATEAREA 0.087 ;
  END WWL

  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9700 1.2000 1.1500 1.4400 ;
        RECT 0.9700 1.0200 1.0650 1.2000 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END RWL

  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0400 1.0950 3.1500 1.4800 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END WBL

  PIN RBL
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0150 0.3500 1.3500 ;
        RECT 0.2500 1.3500 0.4300 1.4400 ;
        RECT 0.2500 0.9200 0.4350 1.0150 ;
        RECT 0.3300 1.4400 0.4300 1.6950 ;
        RECT 0.3350 0.7200 0.4350 0.9200 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END RBL

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 3.1300 1.8050 3.2200 2.0800 ;
        RECT 2.0650 1.3550 2.1550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7250 1.5900 0.9500 1.6850 ;
      RECT 0.7250 1.4200 0.8150 1.5900 ;
      RECT 0.5200 1.3300 0.8800 1.4200 ;
      RECT 0.5200 1.2100 0.6100 1.3300 ;
      RECT 0.7900 0.8750 0.8800 1.3300 ;
      RECT 0.7900 0.7000 0.9250 0.8750 ;
      RECT 0.0700 1.8300 1.4850 1.9200 ;
      RECT 0.0700 0.4800 1.4950 0.5700 ;
      RECT 1.3950 0.5700 1.4950 0.9100 ;
      RECT 0.5950 0.5700 0.6950 0.8900 ;
      RECT 0.0700 1.5000 0.1700 1.8300 ;
      RECT 0.0700 0.8650 0.1600 1.5000 ;
      RECT 0.0700 0.5700 0.1700 0.8650 ;
      RECT 1.8850 1.0750 2.1500 1.2450 ;
      RECT 1.8850 0.7700 2.1050 0.8650 ;
      RECT 1.8850 1.2450 1.9750 1.7950 ;
      RECT 1.8850 0.8650 1.9750 1.0750 ;
      RECT 2.2550 1.8250 2.7000 1.9150 ;
      RECT 2.2550 0.6800 2.3450 1.8250 ;
      RECT 1.6600 0.5900 2.3450 0.6800 ;
      RECT 2.2550 0.5250 2.3450 0.5900 ;
      RECT 2.2550 0.4300 2.5600 0.5250 ;
      RECT 1.6600 0.6800 1.7500 1.0800 ;
      RECT 1.3650 1.0800 1.7500 1.1900 ;
      RECT 2.8600 0.6800 2.9500 1.5150 ;
      RECT 3.4300 1.7150 3.5200 1.9900 ;
      RECT 2.6750 1.6250 3.5200 1.7150 ;
      RECT 3.4300 0.4300 3.5200 1.6250 ;
      RECT 2.4350 0.6500 2.5250 1.2050 ;
      RECT 2.6750 1.3100 2.7650 1.6250 ;
      RECT 2.4350 1.2050 2.7650 1.3100 ;
  END
END RF1R1WS_X1P4M_A12TH

MACRO RF1R1WS_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 1.1000 0.3200 1.2700 0.3600 ;
        RECT 1.6300 0.3200 1.8000 0.3750 ;
        RECT 1.9400 0.3200 2.1100 0.5000 ;
    END
  END VSS

  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9700 1.2000 1.1500 1.4400 ;
        RECT 0.9700 1.0200 1.0650 1.2000 ;
    END
    ANTENNAGATEAREA 0.1452 ;
  END RWL

  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0400 1.0400 3.1500 1.4800 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END WBL

  PIN RBL
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0150 0.3500 1.3500 ;
        RECT 0.2500 1.3500 0.4300 1.4400 ;
        RECT 0.2500 0.9200 0.4350 1.0150 ;
        RECT 0.3400 1.4400 0.4300 1.6950 ;
        RECT 0.3350 0.7200 0.4350 0.9200 ;
    END
    ANTENNADIFFAREA 0.286 ;
  END RBL

  PIN WWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.5800 2.7500 1.1600 ;
        RECT 2.6500 0.4900 3.3400 0.5800 ;
        RECT 3.2500 0.5800 3.3400 0.9800 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END WWL

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 1.0100 2.0100 1.2250 2.0800 ;
        RECT 3.1300 1.8800 3.2200 2.0800 ;
        RECT 2.0750 1.4050 2.1650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7250 1.5950 0.9500 1.6850 ;
      RECT 0.7250 1.4200 0.8150 1.5950 ;
      RECT 0.5200 1.3300 0.8800 1.4200 ;
      RECT 0.5200 1.2100 0.6100 1.3300 ;
      RECT 0.7900 0.9400 0.8800 1.3300 ;
      RECT 0.7900 0.7400 0.9250 0.9400 ;
      RECT 0.0700 1.8300 1.4300 1.9200 ;
      RECT 1.3300 1.5050 1.4300 1.8300 ;
      RECT 0.0700 0.4800 1.4950 0.5700 ;
      RECT 1.3950 0.5700 1.4950 0.9300 ;
      RECT 0.5950 0.5700 0.6950 0.8900 ;
      RECT 0.0700 1.5000 0.1700 1.8300 ;
      RECT 0.0700 0.8650 0.1600 1.5000 ;
      RECT 0.0700 0.5700 0.1700 0.8650 ;
      RECT 1.8950 1.1550 2.1200 1.2450 ;
      RECT 1.9550 1.0750 2.1200 1.1550 ;
      RECT 1.8950 1.2450 1.9850 1.8800 ;
      RECT 1.9550 0.8050 2.0450 1.0750 ;
      RECT 2.2650 1.8750 2.6800 1.9650 ;
      RECT 2.2650 0.6800 2.3550 1.8750 ;
      RECT 1.6600 0.5900 2.3550 0.6800 ;
      RECT 2.2550 0.5250 2.3550 0.5900 ;
      RECT 2.2550 0.4300 2.5600 0.5250 ;
      RECT 1.6600 0.6800 1.7500 1.0800 ;
      RECT 1.3650 1.0800 1.7500 1.1900 ;
      RECT 2.8600 0.6800 2.9500 1.5850 ;
      RECT 3.4300 1.7850 3.5200 1.9900 ;
      RECT 2.6750 1.6950 3.5200 1.7850 ;
      RECT 3.4300 0.5150 3.5200 1.6950 ;
      RECT 2.4450 0.6500 2.5350 1.2550 ;
      RECT 2.6750 1.3600 2.7650 1.6950 ;
      RECT 2.4450 1.2550 2.7650 1.3600 ;
  END
END RF1R1WS_X2M_A12TH

MACRO RF1R2WS_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.3900 0.3200 0.5600 0.5050 ;
        RECT 2.8900 0.3200 3.1000 0.4700 ;
        RECT 3.5200 0.3200 3.7100 0.3700 ;
        RECT 4.6000 0.3200 4.7000 0.7200 ;
    END
  END VSS

  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9850 4.5500 1.4450 ;
    END
    ANTENNAGATEAREA 0.0777 ;
  END RWL

  PIN WBL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9200 2.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0735 ;
  END WBL2

  PIN WWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3750 1.2500 2.0400 1.3500 ;
        RECT 1.3750 1.2000 1.5450 1.2500 ;
        RECT 1.8700 1.2000 2.0400 1.2500 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END WWL2

  PIN WWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1950 1.6500 1.3950 1.8050 ;
        RECT 0.0950 1.8050 1.3950 1.8950 ;
    END
    ANTENNAGATEAREA 0.0774 ;
  END WWL1

  PIN WBL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0050 0.5500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0735 ;
  END WBL1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.3750 2.0100 0.5450 2.0800 ;
        RECT 2.9300 1.9750 3.1000 2.0800 ;
        RECT 3.5650 1.7600 3.6650 2.0800 ;
        RECT 4.6000 1.7000 4.7000 2.0800 ;
    END
  END VDD

  PIN RBL
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0100 1.5900 4.1800 1.7900 ;
        RECT 4.0900 1.7900 4.1800 1.9900 ;
        RECT 4.0100 0.7800 4.1000 1.5900 ;
        RECT 4.0100 0.6900 4.1800 0.7800 ;
        RECT 4.0900 0.4100 4.1800 0.6900 ;
    END
    ANTENNADIFFAREA 0.2288 ;
  END RBL
  OBS
    LAYER M1 ;
      RECT 0.6400 1.4150 0.8100 1.7050 ;
      RECT 0.6400 0.8850 0.7300 1.4150 ;
      RECT 0.6400 0.7950 0.8200 0.8850 ;
      RECT 0.0550 0.5950 1.0000 0.6850 ;
      RECT 0.9100 0.6850 1.0000 1.3300 ;
      RECT 0.0550 1.5000 0.1700 1.7100 ;
      RECT 0.0550 0.8550 0.1450 1.5000 ;
      RECT 0.0550 0.6850 0.1700 0.8550 ;
      RECT 2.1600 1.3200 2.2500 1.6100 ;
      RECT 2.1600 1.1500 2.3250 1.3200 ;
      RECT 2.1600 0.7600 2.2500 1.1500 ;
      RECT 1.4250 0.6700 2.2500 0.7600 ;
      RECT 1.4250 0.7600 1.5150 1.0900 ;
      RECT 2.6100 1.6000 2.8400 1.6900 ;
      RECT 2.6100 0.8300 2.7000 1.6000 ;
      RECT 2.6100 0.7400 2.8250 0.8300 ;
      RECT 1.5850 1.8850 2.8550 1.9200 ;
      RECT 1.5850 1.8300 3.3200 1.8850 ;
      RECT 2.7650 1.7950 3.3200 1.8300 ;
      RECT 3.2300 0.7650 3.3200 1.7950 ;
      RECT 1.5850 1.7950 1.7550 1.8300 ;
      RECT 1.0900 0.5600 3.5350 0.5700 ;
      RECT 2.4150 0.5700 3.5350 0.6500 ;
      RECT 3.4450 0.6500 3.5350 1.0250 ;
      RECT 3.4450 1.0250 3.7350 1.1950 ;
      RECT 1.0900 0.4800 2.5050 0.5600 ;
      RECT 2.4150 0.6500 2.5050 1.7200 ;
      RECT 0.9800 1.4450 1.1800 1.5350 ;
      RECT 1.0900 0.5700 1.1800 1.4450 ;
      RECT 3.8300 0.4950 3.9200 1.9400 ;
      RECT 4.2700 1.7150 4.4700 1.8100 ;
      RECT 4.2700 0.6100 4.4950 0.7000 ;
      RECT 4.2700 1.4800 4.3600 1.7150 ;
      RECT 4.1900 1.3900 4.3600 1.4800 ;
      RECT 4.1900 0.9800 4.2800 1.3900 ;
      RECT 4.1900 0.8900 4.3600 0.9800 ;
      RECT 4.2700 0.7000 4.3600 0.8900 ;
  END
END RF1R2WS_X1M_A12TH

MACRO RF1R2WS_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.4450 ;
        RECT 3.1900 0.3200 3.4000 0.4900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 1.8350 1.7800 1.9350 2.0800 ;
        RECT 2.1400 1.7800 2.2400 2.0800 ;
        RECT 3.2600 1.7000 3.3600 2.0800 ;
    END
  END VDD

  PIN WBL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9650 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END WBL1

  PIN WWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.5750 1.3500 1.4600 ;
        RECT 0.2700 0.5350 1.3500 0.5750 ;
        RECT 0.2700 0.5750 0.9650 0.6250 ;
        RECT 0.8400 0.4850 1.3500 0.5350 ;
        RECT 0.8750 0.6250 0.9650 0.9100 ;
        RECT 0.2700 0.6250 0.3600 0.7300 ;
        RECT 0.8500 0.9100 0.9650 1.0800 ;
        RECT 0.2550 0.7300 0.3600 0.9000 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END WWL1

  PIN WWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 1.0100 2.3650 1.1900 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END WWL2

  PIN WBL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0750 1.2500 3.3900 1.3500 ;
        RECT 3.0750 1.0000 3.1750 1.2500 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END WBL2

  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0100 4.1500 1.4300 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END RWL

  PIN RBL
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4100 1.0500 4.7150 1.1500 ;
        RECT 4.6250 1.1500 4.7150 1.6350 ;
        RECT 4.6250 0.9000 4.7150 1.0500 ;
        RECT 4.5050 1.6350 4.7150 1.7250 ;
        RECT 4.5650 0.8100 4.7150 0.9000 ;
        RECT 4.5650 0.4650 4.6550 0.8100 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END RBL
  OBS
    LAYER M1 ;
      RECT 0.6400 1.3000 0.7450 1.4850 ;
      RECT 0.6400 0.8250 0.7300 1.3000 ;
      RECT 0.5950 0.7350 0.7850 0.8250 ;
      RECT 0.0500 1.6250 0.9650 1.7150 ;
      RECT 0.8750 1.1900 0.9650 1.6250 ;
      RECT 0.0500 1.7150 0.1700 1.8500 ;
      RECT 0.0500 0.6250 0.1400 1.6250 ;
      RECT 0.0500 0.4550 0.1700 0.6250 ;
      RECT 1.8100 1.1300 1.9000 1.4550 ;
      RECT 1.6600 1.0400 1.9000 1.1300 ;
      RECT 1.8100 0.7250 1.9000 1.0400 ;
      RECT 2.4000 1.3500 2.6250 1.4400 ;
      RECT 2.5350 0.9000 2.6250 1.3500 ;
      RECT 2.4600 0.8100 2.6250 0.9000 ;
      RECT 2.4600 0.5750 2.5500 0.8100 ;
      RECT 1.4500 0.4850 2.5500 0.5750 ;
      RECT 1.4500 0.5750 1.5400 0.9000 ;
      RECT 2.8950 0.7750 3.1250 0.8650 ;
      RECT 2.8950 1.4600 3.0650 1.8500 ;
      RECT 2.8950 0.8650 2.9850 1.4600 ;
      RECT 2.7150 0.5800 3.4350 0.6700 ;
      RECT 3.3450 0.6700 3.4350 1.1400 ;
      RECT 1.0550 1.6600 1.1450 1.9500 ;
      RECT 1.0550 0.6850 1.1450 1.5700 ;
      RECT 1.0550 1.5700 2.8050 1.6600 ;
      RECT 2.7150 1.6600 2.8050 1.7400 ;
      RECT 2.7150 0.6700 2.8050 1.5700 ;
      RECT 4.3050 1.3050 4.5350 1.3950 ;
      RECT 3.7350 1.6350 4.3950 1.7250 ;
      RECT 4.3050 1.3950 4.3950 1.6350 ;
      RECT 3.7350 0.6600 4.1950 0.7500 ;
      RECT 3.7350 0.7500 3.8250 1.6350 ;
      RECT 3.5250 1.8150 4.9150 1.9050 ;
      RECT 4.8250 0.4650 4.9150 1.8150 ;
      RECT 3.5250 0.4800 4.3950 0.5700 ;
      RECT 4.3050 0.5700 4.3950 0.8700 ;
      RECT 4.3050 0.4100 4.3950 0.4800 ;
      RECT 3.5250 0.5700 3.6150 1.8150 ;
  END
END RF1R2WS_X1P4M_A12TH

MACRO RF1R2WS_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.4450 ;
        RECT 0.8900 0.3200 1.0600 0.4450 ;
        RECT 3.6500 0.3200 3.8600 0.4900 ;
        RECT 4.2000 0.3200 4.4100 0.4900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 0.3350 1.8750 0.5450 2.0800 ;
        RECT 0.8550 1.8750 1.0650 2.0800 ;
        RECT 2.2650 1.7800 2.3650 2.0800 ;
        RECT 2.6250 1.7800 2.7250 2.0800 ;
        RECT 3.7500 1.7250 3.8500 2.0800 ;
        RECT 4.2700 1.7250 4.3700 2.0800 ;
    END
  END VDD

  PIN WBL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0350 0.5500 1.4600 ;
    END
    ANTENNAGATEAREA 0.1194 ;
  END WBL1

  PIN WWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7450 1.2500 1.9950 1.3500 ;
        RECT 1.7450 0.5750 1.8450 1.2500 ;
        RECT 0.2600 0.5350 1.8450 0.5750 ;
        RECT 0.2600 0.5750 1.4300 0.6250 ;
        RECT 1.2750 0.4850 1.8450 0.5350 ;
        RECT 0.2600 0.6250 0.3500 0.7500 ;
        RECT 1.3400 0.6250 1.4300 1.0400 ;
        RECT 0.2350 0.7500 0.3500 0.9200 ;
        RECT 1.1900 1.0400 1.4300 1.1300 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END WWL1

  PIN WWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0100 2.8500 1.1900 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END WWL2

  PIN WBL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0750 1.2500 4.3900 1.3500 ;
        RECT 4.0750 1.0000 4.1750 1.2500 ;
    END
    ANTENNAGATEAREA 0.1194 ;
  END WBL2

  PIN RWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.0100 5.1500 1.4300 ;
    END
    ANTENNAGATEAREA 0.1194 ;
  END RWL

  PIN RBL
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4100 1.0500 5.7400 1.1500 ;
        RECT 5.6500 1.1500 5.7400 1.6350 ;
        RECT 5.6500 0.8850 5.7400 1.0500 ;
        RECT 5.5100 1.6350 5.7400 1.7250 ;
        RECT 5.5700 0.4650 5.7400 0.8850 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END RBL
  OBS
    LAYER M1 ;
      RECT 0.6550 1.5150 1.2700 1.6050 ;
      RECT 1.1800 1.4100 1.2700 1.5150 ;
      RECT 0.6150 0.8300 1.2500 0.9200 ;
      RECT 1.1600 0.7350 1.2500 0.8300 ;
      RECT 0.6550 0.9200 0.7450 1.5150 ;
      RECT 0.6150 0.7150 0.7850 0.8300 ;
      RECT 0.0500 1.6950 1.4550 1.7850 ;
      RECT 1.3650 1.2200 1.4550 1.6950 ;
      RECT 0.0500 1.7850 0.1700 1.8950 ;
      RECT 0.0500 0.6250 0.1400 1.6950 ;
      RECT 0.0500 0.4550 0.1700 0.6250 ;
      RECT 2.2600 1.3050 2.4500 1.3950 ;
      RECT 2.2600 1.1000 2.3500 1.3050 ;
      RECT 2.1050 1.0100 2.3500 1.1000 ;
      RECT 2.2600 0.8550 2.3500 1.0100 ;
      RECT 2.2600 0.7650 2.4500 0.8550 ;
      RECT 2.8850 1.4000 3.1100 1.4900 ;
      RECT 3.0200 0.8950 3.1100 1.4000 ;
      RECT 2.9450 0.8050 3.1100 0.8950 ;
      RECT 2.9450 0.5850 3.0350 0.8050 ;
      RECT 1.9350 0.4950 3.0350 0.5850 ;
      RECT 1.9350 0.5850 2.0250 0.7000 ;
      RECT 3.4100 1.4400 4.1050 1.5300 ;
      RECT 4.0150 1.5300 4.1050 1.8550 ;
      RECT 3.4100 0.7750 4.1300 0.8650 ;
      RECT 3.4600 1.5300 3.5500 1.8500 ;
      RECT 3.4100 0.8650 3.5000 1.4400 ;
      RECT 3.2000 0.5800 4.4450 0.6700 ;
      RECT 4.3550 0.6700 4.4450 1.1400 ;
      RECT 1.5450 1.6900 1.6350 1.9500 ;
      RECT 1.5650 0.9550 1.6550 1.6000 ;
      RECT 1.5200 0.7450 1.6550 0.9550 ;
      RECT 2.3350 1.5650 2.5050 1.6000 ;
      RECT 1.5450 1.6000 3.2900 1.6900 ;
      RECT 3.2000 1.6900 3.2900 1.8350 ;
      RECT 3.2000 0.6700 3.2900 1.6000 ;
      RECT 5.3100 1.3050 5.5600 1.3950 ;
      RECT 4.7350 1.6500 5.4000 1.7400 ;
      RECT 5.3100 1.3950 5.4000 1.6500 ;
      RECT 4.7350 0.6600 5.2000 0.7500 ;
      RECT 4.7350 0.7500 4.8250 1.6500 ;
      RECT 4.5350 1.8300 5.9200 1.9200 ;
      RECT 5.8300 0.4650 5.9200 1.8300 ;
      RECT 4.5350 0.4800 5.4000 0.5700 ;
      RECT 5.3100 0.5700 5.4000 0.9000 ;
      RECT 4.5350 0.5700 4.6250 1.8300 ;
  END
END RF1R2WS_X2M_A12TH

MACRO RF2R1WS_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3500 0.3200 0.5200 0.4800 ;
        RECT 1.5950 0.3200 1.9650 0.3750 ;
        RECT 2.9150 0.3200 3.0850 0.5750 ;
        RECT 4.0100 0.3200 4.1100 0.8550 ;
    END
  END VSS

  PIN RBL2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.5400 3.5650 0.9700 ;
        RECT 3.4500 0.9700 3.5500 1.4400 ;
        RECT 3.4500 1.4400 3.5650 1.8700 ;
    END
    ANTENNADIFFAREA 0.25025 ;
  END RBL2

  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.1500 2.3500 1.4350 ;
        RECT 2.2500 1.4350 2.4500 1.5350 ;
        RECT 2.2500 1.0500 2.4500 1.1500 ;
        RECT 2.3500 1.5350 2.4500 1.9350 ;
        RECT 2.3500 0.8050 2.4500 1.0500 ;
    END
    ANTENNADIFFAREA 0.239525 ;
  END RBL1

  PIN RWL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1500 4.1500 1.3900 ;
        RECT 3.8800 1.0500 4.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0777 ;
  END RWL2

  PIN RWL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.3350 2.9500 1.6100 ;
        RECT 2.7300 1.2450 2.9500 1.3350 ;
    END
    ANTENNAGATEAREA 0.0777 ;
  END RWL1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 2.9500 1.8400 3.0500 2.0800 ;
        RECT 4.0100 1.6350 4.1100 2.0800 ;
    END
  END VDD

  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0250 0.5800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END WBL

  PIN WWL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8200 0.3500 1.2400 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END WWL
  OBS
    LAYER M1 ;
      RECT 2.5400 0.8500 2.7550 0.9400 ;
      RECT 2.6200 1.5750 2.7100 1.6900 ;
      RECT 2.5400 1.4850 2.7100 1.5750 ;
      RECT 2.5400 0.9400 2.6300 1.4850 ;
      RECT 1.0750 0.6700 3.1250 0.6950 ;
      RECT 2.5850 0.6950 3.1250 0.7600 ;
      RECT 3.0350 0.7600 3.1250 1.2150 ;
      RECT 1.0750 0.6050 2.6750 0.6700 ;
      RECT 0.8900 1.6250 1.9100 1.7150 ;
      RECT 1.8200 0.6950 1.9100 1.6250 ;
      RECT 1.0750 0.5050 1.1650 0.6050 ;
      RECT 0.9450 0.4150 1.1650 0.5050 ;
      RECT 3.2150 0.5400 3.3050 1.8700 ;
      RECT 3.7550 1.6000 3.8450 1.7150 ;
      RECT 3.6600 1.5100 3.8450 1.6000 ;
      RECT 3.6600 0.9400 3.7500 1.5100 ;
      RECT 3.6600 0.8500 3.8450 0.9400 ;
      RECT 3.7550 0.6850 3.8450 0.8500 ;
      RECT 0.6900 0.8050 0.7800 1.7150 ;
      RECT 0.1100 1.8300 1.3100 1.9200 ;
      RECT 0.0500 0.5950 0.9650 0.6850 ;
      RECT 0.8750 0.6850 0.9650 0.8500 ;
      RECT 0.8750 0.8500 1.3100 0.9400 ;
      RECT 0.8750 0.9400 0.9650 1.2900 ;
      RECT 0.8750 1.2900 1.0650 1.3800 ;
      RECT 0.0500 1.3200 0.1700 1.6900 ;
      RECT 0.0500 0.6850 0.1400 1.3200 ;
      RECT 0.0950 0.4100 0.1850 0.5950 ;
      RECT 1.5450 1.1750 1.6350 1.4500 ;
      RECT 1.3500 1.0850 1.6350 1.1750 ;
      RECT 1.5450 0.8050 1.6350 1.0850 ;
      RECT 2.0950 1.6900 2.1850 1.9900 ;
      RECT 2.0100 1.6000 2.1850 1.6900 ;
      RECT 2.0100 0.9350 2.1000 1.6000 ;
      RECT 2.0100 0.8450 2.2450 0.9350 ;
  END
END RF2R1WS_X1M_A12TH

MACRO OR6_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.4750 ;
        RECT 0.9100 0.3200 1.0100 0.4750 ;
        RECT 2.0250 0.3200 2.1250 0.3900 ;
        RECT 2.5850 0.3200 2.6750 0.4750 ;
        RECT 3.1250 0.3200 3.2150 0.4750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.0900 1.6750 0.1900 2.0800 ;
        RECT 1.5000 1.6700 1.6100 2.0800 ;
        RECT 2.0450 1.6700 2.1350 2.0800 ;
        RECT 3.4150 1.6700 3.5250 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 0.8500 1.2000 0.9500 ;
        RECT 1.1000 0.9500 1.2000 1.1400 ;
        RECT 0.4000 0.8250 0.6200 0.8500 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.2500 1.4000 1.3500 ;
        RECT 1.3000 1.2100 1.4000 1.2500 ;
        RECT 0.2000 1.2050 0.3000 1.2500 ;
        RECT 1.3000 1.1100 1.4700 1.2100 ;
        RECT 0.0850 1.1050 0.3000 1.2050 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8000 1.9500 1.3400 ;
        RECT 1.7650 1.3400 1.9500 1.4400 ;
        RECT 1.4700 0.7000 1.9500 0.8000 ;
        RECT 1.7650 1.4400 1.8650 1.7850 ;
        RECT 1.4700 0.6600 1.6400 0.7000 ;
    END
    ANTENNADIFFAREA 0.285 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0500 3.0700 1.1500 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END D

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2200 1.2500 3.4000 1.3500 ;
        RECT 3.3000 1.2100 3.4000 1.2500 ;
        RECT 2.2200 1.0500 2.3200 1.2500 ;
        RECT 3.3000 1.1100 3.5100 1.2100 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END F

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4400 0.8500 3.2000 0.9500 ;
        RECT 2.4400 0.9500 2.5400 1.1250 ;
        RECT 2.9900 0.7950 3.2000 0.8500 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END E
  OBS
    LAYER M1 ;
      RECT 0.7750 1.4850 1.6750 1.5750 ;
      RECT 1.5850 1.0000 1.6750 1.4850 ;
      RECT 1.2900 0.9100 1.6750 1.0000 ;
      RECT 1.2900 0.6950 1.3800 0.9100 ;
      RECT 0.0900 0.6050 1.3800 0.6950 ;
      RECT 0.0900 0.4550 0.1900 0.6000 ;
      RECT 0.7750 1.5750 0.8650 1.9150 ;
      RECT 0.0900 0.6950 0.7500 0.7000 ;
      RECT 0.0900 0.6000 0.7500 0.6050 ;
      RECT 0.6500 0.4550 0.7500 0.6000 ;
      RECT 1.4800 0.5100 2.4600 0.5700 ;
      RECT 1.1950 0.4800 2.4600 0.5100 ;
      RECT 1.1950 0.4200 1.5700 0.4800 ;
      RECT 2.0400 0.6600 3.5150 0.7000 ;
      RECT 2.6000 0.6100 3.5150 0.6600 ;
      RECT 3.4250 0.4550 3.5150 0.6100 ;
      RECT 2.0400 0.7500 2.1300 1.4550 ;
      RECT 2.7850 1.5450 2.8750 1.8850 ;
      RECT 2.0400 1.4550 2.8750 1.5450 ;
      RECT 2.0400 0.7000 2.7000 0.7500 ;
      RECT 2.8650 0.4550 2.9550 0.6100 ;
  END
END OR6_X1P4M_A12TH

MACRO OR6_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 1.1900 0.3200 1.2800 0.5800 ;
        RECT 1.7100 0.3200 1.8000 0.5800 ;
        RECT 2.2300 0.3200 2.3200 0.5600 ;
        RECT 3.3000 0.3200 3.3900 0.5600 ;
        RECT 3.7400 0.3200 3.8300 0.5650 ;
        RECT 4.2900 0.3200 4.3800 0.5650 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 3.7500 1.9900 3.9200 2.0800 ;
        RECT 2.7500 1.8400 2.8400 2.0800 ;
        RECT 1.7100 1.7050 1.8000 2.0800 ;
        RECT 2.2300 1.6200 2.3200 2.0800 ;
        RECT 3.2700 1.6200 3.3600 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1150 1.2500 5.2050 1.3500 ;
    END
    ANTENNAGATEAREA 0.153 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5400 1.2500 3.9600 1.3500 ;
    END
    ANTENNAGATEAREA 0.153 ;
  END C

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7700 1.2300 2.1900 1.3500 ;
    END
    ANTENNAGATEAREA 0.153 ;
  END F

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6250 1.0500 1.4350 1.1500 ;
        RECT 0.6250 1.1500 0.7150 1.2650 ;
        RECT 1.3450 1.1500 1.4350 1.2350 ;
        RECT 1.3350 1.0450 1.4350 1.0500 ;
    END
    ANTENNAGATEAREA 0.153 ;
  END E

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4100 1.0500 4.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.153 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4850 1.4500 3.1000 1.5500 ;
        RECT 2.4850 1.5500 2.5800 1.9800 ;
        RECT 3.0100 1.5500 3.1000 1.9900 ;
        RECT 2.4850 1.0150 2.5750 1.4500 ;
        RECT 2.4850 0.9250 2.8800 1.0150 ;
        RECT 2.7100 0.6650 2.8800 0.9250 ;
    END
    ANTENNADIFFAREA 0.402 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 0.8500 1.0150 0.9500 ;
    END
    ANTENNAGATEAREA 0.153 ;
  END D
  OBS
    LAYER M1 ;
      RECT 1.4450 1.5250 2.0600 1.6150 ;
      RECT 1.9700 1.6150 2.0600 1.9250 ;
      RECT 0.5400 1.9200 0.6300 1.9900 ;
      RECT 0.5400 1.8300 1.5400 1.9200 ;
      RECT 0.5400 1.6200 0.6300 1.8300 ;
      RECT 1.4450 1.6150 1.5400 1.8300 ;
      RECT 2.4550 0.4800 3.1400 0.5700 ;
      RECT 3.0500 0.5700 3.1400 1.0400 ;
      RECT 3.0500 1.0400 3.2450 1.1300 ;
      RECT 2.3050 0.7600 2.3950 1.2800 ;
      RECT 0.8900 0.6700 2.5450 0.7600 ;
      RECT 2.4550 0.5700 2.5450 0.6700 ;
      RECT 0.0800 1.4400 1.0900 1.5300 ;
      RECT 1.0000 1.5300 1.0900 1.7400 ;
      RECT 1.0000 1.4350 1.0900 1.4400 ;
      RECT 0.8900 0.4100 1.0600 0.6700 ;
      RECT 1.0000 1.3450 1.6600 1.4350 ;
      RECT 1.5700 0.7600 1.6600 1.3450 ;
      RECT 1.4100 0.4150 1.5800 0.6700 ;
      RECT 0.0800 1.5300 0.1700 1.9400 ;
      RECT 4.0100 1.9200 4.1800 1.9700 ;
      RECT 4.0100 1.8300 5.1200 1.9200 ;
      RECT 4.0100 1.7450 4.1800 1.8300 ;
      RECT 3.4900 1.6550 4.1800 1.7450 ;
      RECT 3.4900 1.7450 3.6600 1.9700 ;
      RECT 5.4300 1.7400 5.5200 1.8900 ;
      RECT 4.4500 1.6500 5.5200 1.7400 ;
      RECT 5.4300 0.7500 5.5200 1.6500 ;
      RECT 3.3350 0.6600 5.5200 0.7500 ;
      RECT 4.5350 0.4450 4.7050 0.6600 ;
      RECT 3.3350 0.7500 3.4250 1.2550 ;
      RECT 2.7100 1.2550 3.4250 1.3450 ;
      RECT 3.9600 0.4450 4.1300 0.6600 ;
  END
END OR6_X2M_A12TH

MACRO OR6_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.7050 ;
        RECT 0.9250 0.3200 1.0150 0.7050 ;
        RECT 1.5750 0.3200 1.6650 0.7050 ;
        RECT 2.1600 0.3200 2.2500 0.7050 ;
        RECT 3.4850 0.3200 3.5750 0.5600 ;
        RECT 4.0150 0.3200 4.1150 0.6100 ;
        RECT 4.2850 0.3200 4.3750 0.7050 ;
        RECT 4.8700 0.3200 4.9600 0.7050 ;
        RECT 5.5200 0.3200 5.6100 0.7050 ;
        RECT 6.1050 0.3200 6.1950 0.7050 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 1.8950 1.7700 1.9950 2.0800 ;
        RECT 4.5400 1.7700 4.6400 2.0800 ;
        RECT 2.9500 1.5100 3.0500 2.0800 ;
        RECT 3.4850 1.5100 3.5850 2.0800 ;
        RECT 2.4300 1.4800 2.5300 2.0800 ;
        RECT 4.0050 1.4800 4.1050 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0650 1.0500 1.5750 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.0500 0.7350 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7250 1.0500 2.1550 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4300 0.8500 3.3500 0.9500 ;
        RECT 3.2500 0.9500 3.3500 1.3000 ;
        RECT 2.9550 0.7400 3.0450 0.8500 ;
        RECT 2.4300 0.5200 2.5300 0.8500 ;
        RECT 2.6950 1.3000 3.8400 1.3900 ;
        RECT 2.6950 1.3900 2.7850 1.7300 ;
        RECT 3.2150 1.3900 3.3050 1.7300 ;
        RECT 3.7500 1.3900 3.8400 1.7300 ;
    END
    ANTENNADIFFAREA 0.6492 ;
  END Y

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9950 1.0500 5.5050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END E

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8000 1.0500 6.3100 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END D

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2200 1.0500 4.7300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END F
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8300 1.4700 1.9200 ;
      RECT 0.3400 1.5100 0.4300 1.8300 ;
      RECT 0.8600 1.5100 0.9500 1.8300 ;
      RECT 1.3800 1.5100 1.4700 1.8300 ;
      RECT 1.6100 1.5000 2.2500 1.5900 ;
      RECT 2.1600 1.5900 2.2500 1.9400 ;
      RECT 1.6100 1.5900 1.7300 1.9300 ;
      RECT 1.6100 1.3900 1.7000 1.5000 ;
      RECT 1.1200 1.3000 1.7000 1.3900 ;
      RECT 1.1200 1.3900 1.2100 1.7100 ;
      RECT 2.2500 1.0800 3.1100 1.1700 ;
      RECT 0.6000 0.8100 2.3400 0.9000 ;
      RECT 2.2500 0.9000 2.3400 1.0800 ;
      RECT 0.0800 1.3900 0.1700 1.7300 ;
      RECT 0.6000 1.3900 0.6900 1.7100 ;
      RECT 0.6000 0.5100 0.6900 0.8100 ;
      RECT 1.2450 0.5100 1.3350 0.8100 ;
      RECT 0.0800 1.3000 0.9450 1.3900 ;
      RECT 0.8550 0.9000 0.9450 1.3000 ;
      RECT 1.9000 0.5100 1.9900 0.8100 ;
      RECT 3.2150 0.6600 3.8400 0.7500 ;
      RECT 3.7500 0.5400 3.8400 0.6600 ;
      RECT 3.2150 0.5700 3.3050 0.6600 ;
      RECT 2.6350 0.4800 3.3050 0.5700 ;
      RECT 4.2850 1.5000 4.9450 1.5900 ;
      RECT 4.8050 1.5900 4.9450 1.9250 ;
      RECT 4.8550 1.3900 4.9450 1.5000 ;
      RECT 4.8550 1.3000 5.4150 1.3900 ;
      RECT 5.3250 1.3900 5.4150 1.7100 ;
      RECT 4.2850 1.5900 4.3750 1.9300 ;
      RECT 5.0650 1.8300 6.1950 1.9200 ;
      RECT 5.0650 1.5100 5.1550 1.8300 ;
      RECT 5.5850 1.5100 5.6750 1.8300 ;
      RECT 6.1050 1.5100 6.1950 1.8300 ;
      RECT 5.6150 1.3000 6.4550 1.3900 ;
      RECT 6.3650 1.3900 6.4550 1.7300 ;
      RECT 3.9100 0.9000 4.0000 1.0800 ;
      RECT 3.4700 1.0800 4.0000 1.1700 ;
      RECT 4.5450 0.5100 4.6350 0.8100 ;
      RECT 5.2000 0.5100 5.2900 0.8100 ;
      RECT 5.8450 1.3900 5.9350 1.7100 ;
      RECT 3.9100 0.8100 5.9350 0.9000 ;
      RECT 5.8450 0.5100 5.9350 0.8100 ;
      RECT 5.6150 0.9000 5.7050 1.3000 ;
  END
END OR6_X3M_A12TH

MACRO OR6_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.4450 0.3200 ;
        RECT 0.6000 0.3200 0.6900 0.7700 ;
        RECT 1.1200 0.3200 1.2100 0.7500 ;
        RECT 1.9250 0.3200 2.0950 0.4050 ;
        RECT 2.4250 0.3200 2.6350 0.4250 ;
        RECT 3.0050 0.3200 3.0950 0.7300 ;
        RECT 3.2100 0.3200 3.3000 0.3800 ;
        RECT 4.0950 0.3200 4.2650 0.5050 ;
        RECT 5.0600 0.3200 5.1500 0.5600 ;
        RECT 5.3100 0.3200 5.4000 0.6250 ;
        RECT 5.8300 0.3200 5.9200 0.6250 ;
        RECT 6.4300 0.3200 6.6450 0.3700 ;
        RECT 7.1900 0.3200 7.2800 0.7500 ;
        RECT 7.7100 0.3200 7.8000 0.7500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7800 1.4500 4.4500 1.5500 ;
        RECT 4.3600 0.9550 4.4500 1.4500 ;
        RECT 3.7800 0.8900 3.8700 1.4500 ;
        RECT 4.3600 0.8650 4.9100 0.9550 ;
        RECT 3.6050 0.8000 3.8700 0.8900 ;
        RECT 4.8200 0.9550 4.9100 1.5500 ;
    END
    ANTENNADIFFAREA 0.806 ;
  END Y

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 1.0500 0.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END F

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8250 0.5700 6.9500 1.2800 ;
        RECT 6.0100 0.4800 6.9500 0.5700 ;
        RECT 6.0100 0.5700 6.1000 0.8500 ;
        RECT 5.8400 0.8500 6.1000 0.9550 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.5250 1.0500 7.9850 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7450 1.5500 1.1300 ;
        RECT 1.4500 1.1300 1.6600 1.2200 ;
        RECT 1.4500 0.6550 2.0750 0.7450 ;
        RECT 1.9850 0.6050 2.0750 0.6550 ;
        RECT 1.9850 0.5150 2.5550 0.6050 ;
        RECT 2.4650 0.6050 2.5550 1.0500 ;
        RECT 2.4650 1.0500 2.6650 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0500 2.1500 1.6500 ;
        RECT 2.0500 1.6500 3.0950 1.7400 ;
        RECT 3.0050 1.0200 3.0950 1.6500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END E

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 1.3500 6.1500 1.6500 ;
        RECT 5.5600 1.6500 6.1500 1.7400 ;
        RECT 6.0500 1.2600 6.4600 1.3500 ;
        RECT 5.5600 1.3500 5.6500 1.6500 ;
        RECT 6.3700 1.0500 6.4600 1.2600 ;
        RECT 5.4200 1.2600 5.6500 1.3500 ;
        RECT 6.3700 0.8600 6.4750 1.0500 ;
        RECT 5.4200 1.0100 5.5100 1.2600 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.4450 2.7200 ;
        RECT 0.3400 1.8400 0.4300 2.0800 ;
        RECT 0.8600 1.8400 0.9500 2.0800 ;
        RECT 7.4500 1.8400 7.5400 2.0800 ;
        RECT 7.9700 1.8400 8.0600 2.0800 ;
        RECT 3.5200 1.8200 3.6100 2.0800 ;
        RECT 4.0400 1.8200 4.1300 2.0800 ;
        RECT 4.5600 1.8200 4.6500 2.0800 ;
        RECT 5.0800 1.8200 5.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 7.0450 0.8400 7.5400 0.9300 ;
      RECT 7.4500 0.5200 7.5400 0.8400 ;
      RECT 3.5750 1.6400 5.1500 1.7300 ;
      RECT 5.0600 1.4050 5.1500 1.6400 ;
      RECT 5.0600 1.3100 5.3200 1.4050 ;
      RECT 5.2300 0.9000 5.3200 1.3100 ;
      RECT 5.2300 0.8100 5.7500 0.9000 ;
      RECT 5.6600 0.9000 5.7500 1.0800 ;
      RECT 5.5700 0.7000 5.7500 0.8100 ;
      RECT 5.5700 0.4100 5.6600 0.7000 ;
      RECT 6.6450 1.3750 7.1350 1.4650 ;
      RECT 7.0450 0.9300 7.1350 1.3750 ;
      RECT 5.7900 1.1700 5.8800 1.5100 ;
      RECT 6.1900 0.6600 6.7350 0.7500 ;
      RECT 6.6450 0.7500 6.7350 1.3750 ;
      RECT 6.7300 1.4650 6.8200 1.7400 ;
      RECT 5.6600 1.0800 6.2800 1.1700 ;
      RECT 6.1900 0.7500 6.2800 1.0800 ;
      RECT 3.5750 1.0000 3.6650 1.6400 ;
      RECT 4.5800 1.1100 4.6700 1.6400 ;
      RECT 7.1900 1.5500 8.3200 1.6400 ;
      RECT 8.2300 1.6400 8.3200 1.9200 ;
      RECT 5.3300 1.8300 7.2800 1.9200 ;
      RECT 7.1900 1.6400 7.2800 1.8300 ;
      RECT 6.2700 1.5500 6.3600 1.8300 ;
      RECT 5.3300 1.5200 5.4200 1.8300 ;
      RECT 7.7100 1.6400 7.8000 1.9200 ;
      RECT 1.1200 1.8300 3.2750 1.9200 ;
      RECT 3.1850 1.4850 3.2750 1.8300 ;
      RECT 0.0800 1.5500 1.2100 1.6400 ;
      RECT 1.1200 1.6400 1.2100 1.8300 ;
      RECT 0.0800 1.6400 0.1700 1.9400 ;
      RECT 0.6000 1.6400 0.6900 1.9400 ;
      RECT 3.2550 0.6600 5.1200 0.7100 ;
      RECT 3.9600 0.7100 5.1200 0.7500 ;
      RECT 5.0300 0.7500 5.1200 1.2100 ;
      RECT 2.7450 0.8350 3.3450 0.9250 ;
      RECT 3.2550 0.9250 3.3450 1.0400 ;
      RECT 3.2550 0.7100 3.3450 0.8350 ;
      RECT 3.2550 1.0400 3.4050 1.2300 ;
      RECT 0.8600 0.5250 0.9500 0.8400 ;
      RECT 1.2250 0.9300 1.3150 1.3100 ;
      RECT 0.8600 0.8400 1.3150 0.9300 ;
      RECT 1.5800 1.4000 1.6700 1.7200 ;
      RECT 1.2250 1.3100 1.8600 1.4000 ;
      RECT 1.7700 0.9400 1.8600 1.3100 ;
      RECT 2.2450 1.2600 2.8950 1.3500 ;
      RECT 2.5450 1.3500 2.6350 1.4600 ;
      RECT 2.8050 0.9800 2.8950 1.2600 ;
      RECT 2.7450 0.9250 2.8950 0.9800 ;
      RECT 2.7450 0.4550 2.8350 0.8350 ;
      RECT 1.7700 0.8500 2.3550 0.9400 ;
      RECT 2.2450 0.9400 2.3550 1.2600 ;
      RECT 2.1850 0.6950 2.3550 0.8500 ;
      RECT 3.2550 0.6200 4.0500 0.6600 ;
      RECT 3.9600 0.7500 4.0500 1.0750 ;
      RECT 3.9600 1.0750 4.2700 1.1650 ;
  END
END OR6_X4M_A12TH

MACRO OR6_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 14.2450 0.3200 ;
        RECT 0.8600 0.3200 0.9500 0.6900 ;
        RECT 1.3800 0.3200 1.4700 0.6900 ;
        RECT 1.9000 0.3200 1.9900 0.6900 ;
        RECT 2.4200 0.3200 2.5100 0.6900 ;
        RECT 2.9400 0.3200 3.0300 0.6900 ;
        RECT 3.9800 0.3200 4.0700 0.6900 ;
        RECT 4.5000 0.3200 4.5900 0.6900 ;
        RECT 5.0200 0.3200 5.1100 0.6900 ;
        RECT 7.2800 0.3200 7.3700 0.5600 ;
        RECT 7.8000 0.3200 7.8900 0.5600 ;
        RECT 8.3200 0.3200 8.4100 0.5600 ;
        RECT 9.0200 0.3200 9.1100 0.7200 ;
        RECT 9.5400 0.3200 9.6300 0.6900 ;
        RECT 10.0600 0.3200 10.1500 0.6900 ;
        RECT 11.1000 0.3200 11.1900 0.6900 ;
        RECT 11.6200 0.3200 11.7100 0.6900 ;
        RECT 12.1400 0.3200 12.2300 0.6900 ;
        RECT 12.6600 0.3200 12.7500 0.6900 ;
        RECT 13.1800 0.3200 13.2700 0.6900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 14.2450 2.7200 ;
        RECT 6.4950 1.7900 6.5950 2.0800 ;
        RECT 7.0150 1.7900 7.1150 2.0800 ;
        RECT 7.5350 1.7900 7.6350 2.0800 ;
        RECT 8.0550 1.7900 8.1550 2.0800 ;
        RECT 5.9750 1.7700 6.0750 2.0800 ;
        RECT 3.9800 1.7250 4.0700 2.0800 ;
        RECT 4.5000 1.7250 4.5900 2.0800 ;
        RECT 5.0200 1.7250 5.1100 2.0800 ;
        RECT 5.5400 1.7250 5.6400 2.0800 ;
        RECT 8.4800 1.7250 8.5800 2.0800 ;
        RECT 9.0200 1.7250 9.1100 2.0800 ;
        RECT 9.5400 1.7250 9.6300 2.0800 ;
        RECT 10.0600 1.7250 10.1500 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0550 1.0500 3.5450 1.1500 ;
    END
    ANTENNAGATEAREA 0.4623 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 1.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.4623 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8650 1.0500 5.0500 1.1500 ;
    END
    ANTENNAGATEAREA 0.4623 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7150 0.8500 6.9500 0.9500 ;
        RECT 6.8500 0.9500 6.9500 1.4550 ;
        RECT 5.7150 0.7350 5.8150 0.8500 ;
        RECT 6.2000 0.6600 6.3700 0.8500 ;
        RECT 6.7200 0.6600 6.8900 0.8500 ;
        RECT 6.2400 1.4550 7.8900 1.5450 ;
        RECT 6.2400 1.5450 6.3300 1.8850 ;
        RECT 6.7600 1.5450 6.8500 1.8850 ;
        RECT 7.2800 1.5450 7.3700 1.8850 ;
        RECT 7.8000 1.5450 7.8900 1.8850 ;
    END
    ANTENNADIFFAREA 1.19 ;
  END Y

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.7950 1.0500 10.2050 1.1500 ;
    END
    ANTENNAGATEAREA 0.4623 ;
  END F

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.6100 1.0500 13.8900 1.1500 ;
    END
    ANTENNAGATEAREA 0.4623 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.5850 1.0500 12.0750 1.1500 ;
    END
    ANTENNAGATEAREA 0.4623 ;
  END E
  OBS
    LAYER M1 ;
      RECT 7.0200 0.6600 8.7100 0.7500 ;
      RECT 8.5400 0.4600 8.7100 0.6600 ;
      RECT 5.4600 0.4800 7.1100 0.5700 ;
      RECT 7.0200 0.5700 7.1100 0.6600 ;
      RECT 7.5000 0.4600 7.6700 0.6600 ;
      RECT 8.0200 0.4600 8.1900 0.6600 ;
      RECT 5.4600 0.5700 5.5500 0.9100 ;
      RECT 5.9800 0.5700 6.0700 0.6900 ;
      RECT 6.5000 0.5700 6.5900 0.6900 ;
      RECT 8.7600 1.5000 10.4100 1.5900 ;
      RECT 10.3200 1.5900 10.4100 1.9300 ;
      RECT 10.3200 1.3900 10.4100 1.5000 ;
      RECT 10.3200 1.3000 11.9700 1.3900 ;
      RECT 10.8400 1.3900 10.9300 1.7100 ;
      RECT 11.3600 1.3900 11.4500 1.7100 ;
      RECT 11.8800 1.3900 11.9700 1.7100 ;
      RECT 8.7600 1.5900 8.8500 1.9300 ;
      RECT 9.2750 1.5900 9.3750 1.9300 ;
      RECT 9.8000 1.5900 9.8900 1.9300 ;
      RECT 10.5800 1.8300 13.7900 1.9200 ;
      RECT 10.5800 1.5100 10.6700 1.8300 ;
      RECT 11.1000 1.5100 11.1900 1.8300 ;
      RECT 11.6200 1.5100 11.7100 1.8300 ;
      RECT 12.6600 1.5100 12.7500 1.8300 ;
      RECT 13.1800 1.5100 13.2700 1.8300 ;
      RECT 13.7000 1.5100 13.7900 1.8300 ;
      RECT 12.1400 1.4900 12.2300 1.8300 ;
      RECT 12.4000 1.3000 14.0500 1.3900 ;
      RECT 13.4400 1.3900 13.5300 1.7100 ;
      RECT 13.9600 1.3900 14.0500 1.7300 ;
      RECT 8.2550 0.8550 13.5300 0.9000 ;
      RECT 9.2800 0.8100 13.5300 0.8550 ;
      RECT 13.4400 0.6300 13.5300 0.8100 ;
      RECT 8.2550 0.9450 8.3450 1.0800 ;
      RECT 7.2750 1.0800 8.3450 1.1700 ;
      RECT 8.2550 0.9000 9.3700 0.9450 ;
      RECT 9.2800 0.6300 9.3700 0.8100 ;
      RECT 9.8000 0.6300 9.8900 0.8100 ;
      RECT 10.8400 0.6300 10.9300 0.8100 ;
      RECT 10.3200 0.6300 10.4100 0.8100 ;
      RECT 11.3600 0.6300 11.4500 0.8100 ;
      RECT 11.8800 0.6300 11.9700 0.8100 ;
      RECT 12.4000 1.3900 12.4900 1.7100 ;
      RECT 12.4000 0.9000 12.4900 1.3000 ;
      RECT 12.4000 0.6300 12.4900 0.8100 ;
      RECT 12.9200 1.3900 13.0100 1.7100 ;
      RECT 12.9200 0.6300 13.0100 0.8100 ;
      RECT 0.3400 1.8300 3.5500 1.9200 ;
      RECT 0.3400 1.5100 0.4300 1.8300 ;
      RECT 0.8600 1.5100 0.9500 1.8300 ;
      RECT 1.3800 1.5100 1.4700 1.8300 ;
      RECT 2.4200 1.5100 2.5100 1.8300 ;
      RECT 2.9400 1.5100 3.0300 1.8300 ;
      RECT 3.4600 1.5100 3.5500 1.8300 ;
      RECT 1.9000 1.4900 1.9900 1.8300 ;
      RECT 3.7200 1.5000 5.3700 1.5900 ;
      RECT 5.2800 1.5900 5.3700 1.9300 ;
      RECT 3.7200 1.5900 3.8100 1.9150 ;
      RECT 3.7200 1.3900 3.8100 1.5000 ;
      RECT 2.1600 1.3000 3.8100 1.3900 ;
      RECT 2.1600 1.3900 2.2500 1.7100 ;
      RECT 2.6800 1.3900 2.7700 1.7100 ;
      RECT 3.2000 1.3900 3.2900 1.7100 ;
      RECT 4.2400 1.5900 4.3300 1.9300 ;
      RECT 4.7550 1.5900 4.8550 1.9300 ;
      RECT 5.2550 1.0800 6.6700 1.1700 ;
      RECT 0.6000 0.8100 5.3450 0.9000 ;
      RECT 5.2550 0.9000 5.3450 1.0800 ;
      RECT 4.2400 0.6300 4.3300 0.8100 ;
      RECT 4.7600 0.6300 4.8500 0.8100 ;
      RECT 2.1600 0.6300 2.2500 0.8100 ;
      RECT 2.6800 0.6300 2.7700 0.8100 ;
      RECT 3.2000 0.6300 3.2900 0.8100 ;
      RECT 3.7200 0.6300 3.8100 0.8100 ;
      RECT 0.6000 1.3900 0.6900 1.7100 ;
      RECT 0.6000 0.6300 0.6900 0.8100 ;
      RECT 1.1200 1.3900 1.2100 1.7100 ;
      RECT 1.1200 0.6300 1.2100 0.8100 ;
      RECT 0.0800 1.3000 1.7300 1.3900 ;
      RECT 1.6400 1.3900 1.7300 1.7100 ;
      RECT 1.6400 0.9000 1.7300 1.3000 ;
      RECT 1.6400 0.6300 1.7300 0.8100 ;
      RECT 0.0800 1.3900 0.1700 1.7300 ;
  END
END OR6_X6M_A12TH

MACRO POSTICG_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.5750 ;
        RECT 1.4950 0.3200 1.5850 0.7250 ;
        RECT 2.6400 0.3200 2.8500 0.3900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9750 1.2500 2.3150 1.3500 ;
        RECT 2.2250 1.3500 2.3150 1.8300 ;
        RECT 1.9750 0.8650 2.0650 1.2500 ;
        RECT 0.9400 1.8300 2.6750 1.9200 ;
        RECT 0.9400 1.5300 1.0300 1.8300 ;
        RECT 2.5850 1.4000 2.6750 1.8300 ;
        RECT 0.8050 1.4400 1.0300 1.5300 ;
        RECT 2.5850 1.3000 2.9400 1.4000 ;
        RECT 2.8500 1.1850 2.9400 1.3000 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6050 0.8500 2.9150 0.9900 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2300 1.0450 1.6300 1.1500 ;
    END
    ANTENNAGATEAREA 0.0222 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6450 0.1500 1.3500 ;
        RECT 0.0500 1.3500 0.1750 1.4400 ;
        RECT 0.0500 0.5550 0.1700 0.6450 ;
        RECT 0.0750 1.4400 0.1750 1.7200 ;
        RECT 0.0800 0.4100 0.1700 0.5550 ;
    END
    ANTENNADIFFAREA 0.1088 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.8650 2.0100 1.0750 2.0800 ;
        RECT 1.4750 2.0100 1.6850 2.0800 ;
        RECT 0.3400 1.6050 0.4300 2.0800 ;
        RECT 2.7650 1.5900 2.8550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6700 0.4550 0.9550 0.5450 ;
      RECT 0.6250 1.2300 0.7150 1.8000 ;
      RECT 0.2400 1.1400 0.7150 1.2300 ;
      RECT 0.2400 1.0200 0.3500 1.1400 ;
      RECT 0.2600 0.7550 0.3500 1.0200 ;
      RECT 0.2600 0.6650 0.7600 0.7550 ;
      RECT 0.6700 0.5450 0.7600 0.6650 ;
      RECT 0.8500 1.2400 1.6800 1.3300 ;
      RECT 1.5900 1.3300 1.6800 1.4850 ;
      RECT 1.1750 1.6500 1.4050 1.7400 ;
      RECT 1.3150 1.3300 1.4050 1.6500 ;
      RECT 0.8500 0.9350 0.9400 1.2400 ;
      RECT 0.4700 0.8450 0.9400 0.9350 ;
      RECT 0.8500 0.7250 0.9400 0.8450 ;
      RECT 0.8500 0.6350 1.1850 0.7250 ;
      RECT 0.4700 0.9350 0.5600 1.0500 ;
      RECT 2.0450 1.5900 2.1350 1.7200 ;
      RECT 1.7750 1.5000 2.1350 1.5900 ;
      RECT 1.7750 0.6550 2.1750 0.7450 ;
      RECT 1.7750 0.9050 1.8650 1.5000 ;
      RECT 1.0300 0.8150 1.8650 0.9050 ;
      RECT 1.7750 0.7450 1.8650 0.8150 ;
      RECT 1.0300 0.9050 1.1200 1.0250 ;
      RECT 2.4050 0.7500 2.4950 1.7200 ;
      RECT 2.2850 0.6600 2.4950 0.7500 ;
      RECT 3.0300 0.5700 3.1200 1.7750 ;
      RECT 2.2250 0.4800 3.1200 0.5700 ;
      RECT 2.2250 0.4200 2.3950 0.4800 ;
  END
END POSTICG_X0P5B_A12TH

MACRO POSTICG_X0P6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.5900 ;
        RECT 1.4700 0.3200 1.6400 0.6800 ;
        RECT 2.6400 0.3200 2.8500 0.3900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.5100 0.9500 1.7750 ;
        RECT 0.8500 1.7750 2.6800 1.8750 ;
        RECT 0.7100 1.4200 0.9500 1.5100 ;
        RECT 2.2300 1.4250 2.3200 1.7750 ;
        RECT 2.5900 1.4000 2.6800 1.7750 ;
        RECT 0.7100 1.1950 0.8000 1.4200 ;
        RECT 2.0550 1.3350 2.3200 1.4250 ;
        RECT 2.5900 1.3000 2.9400 1.4000 ;
        RECT 2.0550 1.0150 2.1450 1.3350 ;
        RECT 2.8500 1.1000 2.9400 1.3000 ;
        RECT 1.9000 0.9250 2.1450 1.0150 ;
    END
    ANTENNAGATEAREA 0.0675 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6000 0.8700 2.7500 1.1000 ;
        RECT 2.6500 0.6950 2.7500 0.8700 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1650 1.0500 1.5000 1.1500 ;
        RECT 1.3900 0.9700 1.5000 1.0500 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6400 0.1500 1.5550 ;
        RECT 0.0500 1.5550 0.1750 1.6650 ;
        RECT 0.0500 0.5700 0.1750 0.6400 ;
        RECT 0.0750 1.6650 0.1750 1.9850 ;
        RECT 0.0750 0.4200 0.1750 0.5700 ;
    END
    ANTENNADIFFAREA 0.1528 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3400 1.9900 0.4300 2.0800 ;
        RECT 0.8350 1.9650 1.0450 2.0800 ;
        RECT 1.4500 1.9650 1.6600 2.0800 ;
        RECT 2.7700 1.5100 2.8600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7100 0.4300 0.9350 0.5200 ;
      RECT 0.5300 1.3450 0.6200 1.6000 ;
      RECT 0.2400 1.2550 0.6200 1.3450 ;
      RECT 0.2400 1.0400 0.3500 1.2550 ;
      RECT 0.2600 0.7700 0.3500 1.0400 ;
      RECT 0.5300 1.6000 0.7400 1.6900 ;
      RECT 0.2600 0.6800 0.8000 0.7700 ;
      RECT 0.7100 0.5200 0.8000 0.6800 ;
      RECT 1.2000 1.3300 1.7100 1.4000 ;
      RECT 0.8900 1.3100 1.7100 1.3300 ;
      RECT 0.8900 0.9500 0.9800 1.2400 ;
      RECT 0.4700 0.8600 0.9800 0.9500 ;
      RECT 0.8900 0.7000 0.9800 0.8600 ;
      RECT 0.8900 0.6100 1.1350 0.7000 ;
      RECT 1.0450 0.5100 1.1350 0.6100 ;
      RECT 1.2000 1.4000 1.2900 1.6850 ;
      RECT 0.8900 1.2400 1.2900 1.3100 ;
      RECT 0.4700 0.9500 0.5600 1.0700 ;
      RECT 2.0300 1.6050 2.1200 1.6850 ;
      RECT 1.8000 1.5150 2.1200 1.6050 ;
      RECT 1.1250 0.7900 2.0800 0.8350 ;
      RECT 1.7100 0.7450 2.0800 0.7900 ;
      RECT 1.9900 0.5550 2.0800 0.7450 ;
      RECT 1.8000 1.1950 1.8900 1.5150 ;
      RECT 1.7000 1.1050 1.8900 1.1950 ;
      RECT 1.7000 0.8800 1.7900 1.1050 ;
      RECT 1.1250 0.8350 1.7900 0.8800 ;
      RECT 1.1250 0.8800 1.2150 0.9600 ;
      RECT 2.4100 0.7500 2.5000 1.6650 ;
      RECT 2.3300 0.6600 2.5000 0.7500 ;
      RECT 3.0300 0.5700 3.1200 1.7200 ;
      RECT 2.2000 0.4800 3.1200 0.5700 ;
      RECT 2.2000 0.4100 2.3750 0.4800 ;
  END
END POSTICG_X0P6B_A12TH

MACRO POSTICG_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6050 ;
        RECT 1.5250 0.3200 1.6150 0.7000 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.5100 0.9500 1.8250 ;
        RECT 0.8400 1.8250 2.7500 1.9150 ;
        RECT 0.8400 1.4200 1.0300 1.5100 ;
        RECT 2.6500 1.4400 2.7500 1.8250 ;
        RECT 2.2500 1.3850 2.3400 1.8250 ;
        RECT 2.6500 1.3300 2.9400 1.4400 ;
        RECT 2.1100 1.2950 2.3400 1.3850 ;
        RECT 2.1100 0.9700 2.2000 1.2950 ;
        RECT 1.9800 0.8800 2.2000 0.9700 ;
    END
    ANTENNAGATEAREA 0.0705 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.6850 2.7500 1.1600 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3400 1.0500 1.6800 1.1500 ;
        RECT 1.3400 1.0000 1.5500 1.0500 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7800 0.1500 1.5650 ;
        RECT 0.0500 1.5650 0.1750 1.7950 ;
        RECT 0.0500 0.6900 0.1900 0.7800 ;
        RECT 0.0900 0.5050 0.1900 0.6900 ;
    END
    ANTENNADIFFAREA 0.1576 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.8900 2.0050 1.1000 2.0800 ;
        RECT 1.4800 2.0050 1.6900 2.0800 ;
        RECT 2.6600 2.0050 2.8700 2.0800 ;
        RECT 0.4150 1.9250 0.5050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6550 0.4300 0.9850 0.5200 ;
      RECT 0.6600 1.6900 0.7500 1.8100 ;
      RECT 0.6050 1.6000 0.7500 1.6900 ;
      RECT 0.6050 1.3750 0.6950 1.6000 ;
      RECT 0.2500 1.2850 0.6950 1.3750 ;
      RECT 0.2500 1.1650 0.3650 1.2850 ;
      RECT 0.2750 0.9350 0.3650 1.1650 ;
      RECT 0.2750 0.8450 0.7450 0.9350 ;
      RECT 0.6550 0.5200 0.7450 0.8450 ;
      RECT 1.2450 1.3700 1.8200 1.4600 ;
      RECT 1.2450 1.4600 1.3350 1.7350 ;
      RECT 1.2450 1.3300 1.3350 1.3700 ;
      RECT 0.9600 1.2400 1.3350 1.3300 ;
      RECT 0.9600 1.1150 1.0500 1.2400 ;
      RECT 0.4900 1.0250 1.0500 1.1150 ;
      RECT 0.9600 0.7000 1.0500 1.0250 ;
      RECT 0.9600 0.6100 1.2150 0.7000 ;
      RECT 0.4900 1.1150 0.5800 1.1950 ;
      RECT 2.0700 1.6350 2.1600 1.7150 ;
      RECT 1.9300 1.5450 2.1600 1.6350 ;
      RECT 1.7900 0.6350 2.2200 0.7250 ;
      RECT 1.7900 0.8800 1.8800 1.1900 ;
      RECT 1.1600 0.7900 1.8800 0.8800 ;
      RECT 1.7900 0.7250 1.8800 0.7900 ;
      RECT 1.9300 1.2800 2.0200 1.5450 ;
      RECT 1.7900 1.1900 2.0200 1.2800 ;
      RECT 1.1600 0.8800 1.2500 1.0300 ;
      RECT 2.4300 0.7500 2.5200 1.7150 ;
      RECT 2.3300 0.6600 2.5200 0.7500 ;
      RECT 3.0300 0.5700 3.1200 1.7700 ;
      RECT 2.3350 0.5100 3.1200 0.5700 ;
      RECT 2.1350 0.4800 3.1200 0.5100 ;
      RECT 2.1350 0.4100 2.4250 0.4800 ;
  END
END POSTICG_X0P7B_A12TH

MACRO POSTICG_X0P8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7550 ;
        RECT 1.5250 0.3200 1.6150 0.6950 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.5100 0.9500 1.8250 ;
        RECT 0.8400 1.8250 2.7500 1.9150 ;
        RECT 0.8400 1.4200 1.0300 1.5100 ;
        RECT 2.6500 1.4400 2.7500 1.8250 ;
        RECT 2.2500 1.3850 2.3400 1.8250 ;
        RECT 2.6500 1.3300 2.9400 1.4400 ;
        RECT 2.1100 1.2950 2.3400 1.3850 ;
        RECT 2.1100 0.9700 2.2000 1.2950 ;
        RECT 1.9800 0.8800 2.2000 0.9700 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.6850 2.7500 1.1600 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3400 1.0500 1.6800 1.1500 ;
        RECT 1.3400 1.0000 1.5500 1.0500 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7800 0.1500 1.4700 ;
        RECT 0.0500 1.4700 0.1750 1.8800 ;
        RECT 0.0500 0.6900 0.1900 0.7800 ;
        RECT 0.0900 0.4100 0.1900 0.6900 ;
    END
    ANTENNADIFFAREA 0.1798 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.9500 2.0050 1.0400 2.0800 ;
        RECT 1.4800 2.0050 1.6900 2.0800 ;
        RECT 2.6800 2.0050 2.8500 2.0800 ;
        RECT 0.4150 1.9250 0.5050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6550 0.4300 0.9850 0.5200 ;
      RECT 0.6600 1.6900 0.7500 1.8100 ;
      RECT 0.6050 1.6000 0.7500 1.6900 ;
      RECT 0.6050 1.3750 0.6950 1.6000 ;
      RECT 0.2500 1.2850 0.6950 1.3750 ;
      RECT 0.2500 1.1650 0.3650 1.2850 ;
      RECT 0.2750 0.9350 0.3650 1.1650 ;
      RECT 0.2750 0.8450 0.7450 0.9350 ;
      RECT 0.6550 0.5200 0.7450 0.8450 ;
      RECT 1.2450 1.3700 1.8200 1.4600 ;
      RECT 1.2450 1.4600 1.3350 1.7350 ;
      RECT 1.2450 1.3300 1.3350 1.3700 ;
      RECT 0.9600 1.2400 1.3350 1.3300 ;
      RECT 0.9600 1.1150 1.0500 1.2400 ;
      RECT 0.4900 1.0250 1.0500 1.1150 ;
      RECT 0.9600 0.7000 1.0500 1.0250 ;
      RECT 0.9600 0.6100 1.2150 0.7000 ;
      RECT 0.4900 1.1150 0.5800 1.1950 ;
      RECT 2.0700 1.6350 2.1600 1.7150 ;
      RECT 1.9300 1.5450 2.1600 1.6350 ;
      RECT 1.7900 0.6350 2.2200 0.7250 ;
      RECT 1.7900 0.8800 1.8800 1.1900 ;
      RECT 1.1600 0.7900 1.8800 0.8800 ;
      RECT 1.7900 0.7250 1.8800 0.7900 ;
      RECT 1.9300 1.2800 2.0200 1.5450 ;
      RECT 1.7900 1.1900 2.0200 1.2800 ;
      RECT 1.1600 0.8800 1.2500 1.0300 ;
      RECT 2.4300 0.7500 2.5200 1.7150 ;
      RECT 2.3300 0.6600 2.5200 0.7500 ;
      RECT 3.0300 0.5700 3.1200 1.7700 ;
      RECT 2.3350 0.5100 3.1200 0.5700 ;
      RECT 2.1350 0.4800 3.1200 0.5100 ;
      RECT 2.1350 0.4100 2.4250 0.4800 ;
  END
END POSTICG_X0P8B_A12TH

MACRO POSTICG_X11B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6350 ;
        RECT 0.8750 0.3200 0.9650 0.6350 ;
        RECT 1.3950 0.3200 1.4850 0.6350 ;
        RECT 1.9150 0.3200 2.0050 0.6350 ;
        RECT 3.7250 0.3200 3.8150 0.6050 ;
        RECT 4.2450 0.3200 4.3350 0.6050 ;
        RECT 4.7650 0.3200 4.8550 0.7200 ;
        RECT 5.3750 0.3200 5.5450 0.8500 ;
        RECT 6.4350 0.3200 6.5250 0.6350 ;
        RECT 7.9100 0.3200 8.0000 0.6750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 1.1650 6.7500 1.8300 ;
        RECT 4.7150 1.8300 7.7400 1.9200 ;
        RECT 6.5250 1.0750 6.7500 1.1650 ;
        RECT 7.6500 1.3450 7.7400 1.8300 ;
        RECT 4.7150 1.2300 4.8050 1.8300 ;
        RECT 3.6600 1.1400 4.8050 1.2300 ;
    END
    ANTENNAGATEAREA 0.4077 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0500 1.0100 8.1750 1.3600 ;
    END
    ANTENNAGATEAREA 0.0885 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1900 1.2500 5.7050 1.3500 ;
    END
    ANTENNAGATEAREA 0.102 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4200 0.9150 0.5800 1.4200 ;
        RECT 0.0950 1.4200 2.7850 1.5800 ;
        RECT 0.0950 0.7550 1.7450 0.9150 ;
        RECT 0.0950 1.5800 0.1850 1.8500 ;
        RECT 0.6150 1.5800 0.7050 1.8500 ;
        RECT 1.1350 1.5800 1.2250 1.8500 ;
        RECT 1.6550 1.5800 1.7450 1.8500 ;
        RECT 2.1750 1.5800 2.2650 1.8500 ;
        RECT 2.6950 1.5800 2.7850 1.8500 ;
        RECT 0.0950 0.4850 0.1850 0.7550 ;
        RECT 0.6150 0.4850 0.7050 0.7550 ;
        RECT 1.1350 0.4850 1.2250 0.7550 ;
        RECT 1.6550 0.4850 1.7450 0.7550 ;
    END
    ANTENNADIFFAREA 1.638875 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.4450 2.7200 ;
        RECT 4.5700 2.0100 4.9800 2.0800 ;
        RECT 5.4100 2.0100 5.5800 2.0800 ;
        RECT 6.0050 2.0100 6.3750 2.0800 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
        RECT 1.9150 1.7700 2.0050 2.0800 ;
        RECT 2.4350 1.7700 2.5250 2.0800 ;
        RECT 3.0500 1.7700 3.1400 2.0800 ;
        RECT 7.8500 1.7700 7.9400 2.0800 ;
        RECT 3.6750 1.6550 3.8450 2.0800 ;
        RECT 4.1950 1.6550 4.3650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.2650 1.3800 4.5850 1.4700 ;
      RECT 4.4950 1.4700 4.5850 1.8400 ;
      RECT 2.1650 0.5400 2.2550 0.6600 ;
      RECT 3.4550 1.4700 3.5450 1.8500 ;
      RECT 3.2650 1.1400 3.3550 1.3800 ;
      RECT 1.2250 1.0500 3.3550 1.1400 ;
      RECT 3.2650 0.7500 3.3550 1.0500 ;
      RECT 2.1650 0.6600 3.3550 0.7500 ;
      RECT 3.9750 1.4700 4.0650 1.8400 ;
      RECT 3.4650 0.7100 4.5950 0.8000 ;
      RECT 4.5050 0.5150 4.5950 0.7100 ;
      RECT 3.4650 0.5700 3.5550 0.7100 ;
      RECT 2.3650 0.4800 3.5550 0.5700 ;
      RECT 3.9850 0.5150 4.0750 0.7100 ;
      RECT 5.1550 0.9400 5.7650 1.0300 ;
      RECT 5.6750 0.6200 5.7650 0.9400 ;
      RECT 5.6750 0.5300 6.2850 0.6200 ;
      RECT 6.1950 0.6200 6.2850 0.7550 ;
      RECT 5.1550 0.5500 5.2450 0.9400 ;
      RECT 4.9150 1.6500 6.0250 1.7400 ;
      RECT 5.9350 1.5300 6.0250 1.6500 ;
      RECT 5.9350 1.4400 6.4350 1.5300 ;
      RECT 6.3450 1.2750 6.4350 1.4400 ;
      RECT 5.9350 0.7600 6.0250 1.4400 ;
      RECT 4.9150 0.9800 5.0050 1.6500 ;
      RECT 4.0250 0.8900 5.0050 0.9800 ;
      RECT 6.1150 0.8450 7.0650 0.9350 ;
      RECT 6.8700 0.9350 6.9600 1.6150 ;
      RECT 6.9750 0.4500 7.0650 0.8450 ;
      RECT 6.1150 0.9350 6.2050 1.2600 ;
      RECT 7.3700 1.6500 7.5400 1.7400 ;
      RECT 7.4500 1.0250 7.5400 1.6500 ;
      RECT 7.4500 0.9350 7.6200 1.0250 ;
      RECT 7.5300 0.6800 7.6200 0.9350 ;
      RECT 8.1700 1.5900 8.2600 1.9350 ;
      RECT 7.8300 1.5000 8.2600 1.5900 ;
      RECT 7.7100 0.8050 8.2600 0.8950 ;
      RECT 8.1700 0.4300 8.2600 0.8050 ;
      RECT 7.8300 0.8950 7.9200 1.5000 ;
      RECT 7.7100 0.5700 7.8000 0.8050 ;
      RECT 7.2350 0.4800 7.8000 0.5700 ;
      RECT 7.2350 0.5700 7.3250 1.0100 ;
      RECT 7.1700 1.0100 7.3250 1.1000 ;
      RECT 7.1700 1.1000 7.2600 1.4050 ;
      RECT 7.0900 1.4050 7.2600 1.7250 ;
  END
END POSTICG_X11B_A12TH

MACRO POSTICG_X13B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 9.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6600 ;
        RECT 0.8750 0.3200 0.9650 0.6600 ;
        RECT 1.3950 0.3200 1.4850 0.6600 ;
        RECT 1.9150 0.3200 2.0050 0.6600 ;
        RECT 4.2600 0.3200 4.3500 0.7100 ;
        RECT 4.7800 0.3200 4.8700 0.7550 ;
        RECT 5.3000 0.3200 5.3900 0.7550 ;
        RECT 6.2500 0.3200 6.3400 0.8800 ;
        RECT 7.2650 0.3200 7.3550 0.6500 ;
        RECT 8.7100 0.3200 8.8000 0.7200 ;
        RECT 9.2300 0.3200 9.3200 0.9000 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4100 1.2500 5.5850 1.3500 ;
        RECT 5.4950 1.3500 5.5850 1.8300 ;
        RECT 4.4100 1.3500 5.1000 1.3650 ;
        RECT 5.4950 1.8300 8.6000 1.9200 ;
        RECT 7.3950 1.8200 8.6000 1.8300 ;
        RECT 7.3950 1.2150 7.4850 1.8200 ;
        RECT 8.5100 1.0500 8.6000 1.8200 ;
        RECT 7.3950 1.1250 7.6050 1.2150 ;
    END
    ANTENNAGATEAREA 0.495 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.8900 1.0400 9.3050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0100 1.2050 6.3800 1.3050 ;
        RECT 6.0100 1.3050 6.1900 1.3500 ;
    END
    ANTENNAGATEAREA 0.12 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 0.9900 0.7900 1.4100 ;
        RECT 0.0950 1.4100 3.3050 1.5900 ;
        RECT 0.0950 0.8100 2.2650 0.9900 ;
        RECT 0.0950 1.5900 0.1850 1.8400 ;
        RECT 0.6150 1.5900 0.7050 1.8400 ;
        RECT 1.1350 1.5900 1.2250 1.8400 ;
        RECT 1.6550 1.5900 1.7450 1.8400 ;
        RECT 2.1750 1.5900 2.2650 1.8400 ;
        RECT 2.6950 1.5900 2.7850 1.8400 ;
        RECT 3.2150 1.5900 3.3050 1.8400 ;
        RECT 0.0950 0.5400 0.1850 0.8100 ;
        RECT 0.6150 0.5400 0.7050 0.8100 ;
        RECT 1.1350 0.5400 1.2250 0.8100 ;
        RECT 1.6550 0.5400 1.7450 0.8100 ;
        RECT 2.1750 0.5350 2.2650 0.8100 ;
    END
    ANTENNADIFFAREA 1.94235 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 9.4450 2.7200 ;
        RECT 6.2350 2.0100 6.4050 2.0800 ;
        RECT 6.7550 2.0100 7.1250 2.0800 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
        RECT 1.9150 1.7700 2.0050 2.0800 ;
        RECT 2.4350 1.7700 2.5250 2.0800 ;
        RECT 2.9550 1.7700 3.0450 2.0800 ;
        RECT 3.4750 1.7700 3.5650 2.0800 ;
        RECT 3.9750 1.6950 4.1450 2.0800 ;
        RECT 4.4950 1.6950 4.6650 2.0800 ;
        RECT 5.0150 1.6950 5.1850 2.0800 ;
        RECT 8.7100 1.4700 8.8000 2.0800 ;
        RECT 9.2300 1.4000 9.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.7550 1.5000 5.4050 1.5900 ;
      RECT 5.3150 1.5900 5.4050 1.9300 ;
      RECT 2.7000 0.6600 2.7900 0.8600 ;
      RECT 3.2300 0.9500 3.3200 1.1300 ;
      RECT 3.2200 0.6600 3.3100 0.8600 ;
      RECT 3.7550 1.5900 3.8450 1.9400 ;
      RECT 3.7550 1.2200 3.8450 1.5000 ;
      RECT 1.2400 1.1300 3.8450 1.2200 ;
      RECT 2.7000 0.8600 3.8300 0.9500 ;
      RECT 3.7400 0.6600 3.8300 0.8600 ;
      RECT 4.2750 1.5900 4.3650 1.9300 ;
      RECT 4.7950 1.5900 4.8850 1.9300 ;
      RECT 4.0000 0.8450 5.6500 0.9350 ;
      RECT 5.5600 0.4350 5.6500 0.8450 ;
      RECT 4.0000 0.5700 4.0900 0.8450 ;
      RECT 2.3800 0.4800 4.0900 0.5700 ;
      RECT 2.9200 0.5700 3.0900 0.7700 ;
      RECT 3.4400 0.5700 3.6100 0.7700 ;
      RECT 4.5200 0.4600 4.6100 0.8450 ;
      RECT 5.0400 0.4600 5.1300 0.8450 ;
      RECT 5.9500 0.9700 6.6350 1.0600 ;
      RECT 6.5450 0.5700 6.6350 0.9700 ;
      RECT 6.5450 0.4800 7.0950 0.5700 ;
      RECT 7.0050 0.5700 7.0950 0.7450 ;
      RECT 7.0050 0.7450 7.2150 0.8350 ;
      RECT 5.9500 0.5400 6.0400 0.9700 ;
      RECT 5.6950 1.6400 6.8350 1.7300 ;
      RECT 6.7450 1.5550 6.8350 1.6400 ;
      RECT 6.7450 1.4650 7.2850 1.5550 ;
      RECT 7.1950 1.3450 7.2850 1.4650 ;
      RECT 6.7450 0.8600 6.8350 1.4650 ;
      RECT 6.7450 0.7700 6.8950 0.8600 ;
      RECT 6.8050 0.6600 6.8950 0.7700 ;
      RECT 5.6950 1.1200 5.7850 1.6400 ;
      RECT 4.6450 1.0300 5.7850 1.1200 ;
      RECT 7.2150 0.9250 7.8400 1.0150 ;
      RECT 7.7500 1.0150 7.8400 1.6650 ;
      RECT 7.7500 0.4400 7.8400 0.9250 ;
      RECT 6.9600 1.0500 7.3050 1.1400 ;
      RECT 7.2150 1.0150 7.3050 1.0500 ;
      RECT 6.9600 1.1400 7.0500 1.2600 ;
      RECT 8.3300 1.1750 8.4200 1.7000 ;
      RECT 8.2600 0.9650 8.4200 1.1750 ;
      RECT 8.3300 0.6950 8.4200 0.9650 ;
      RECT 8.9700 1.3800 9.0600 1.7700 ;
      RECT 8.6900 1.2900 9.0600 1.3800 ;
      RECT 8.5100 0.8100 9.0600 0.9000 ;
      RECT 8.9700 0.4650 9.0600 0.8100 ;
      RECT 8.6900 0.9000 8.7800 1.2900 ;
      RECT 8.5100 0.5700 8.6000 0.8100 ;
      RECT 8.0400 0.4800 8.6000 0.5700 ;
      RECT 8.0400 0.5700 8.1300 0.8600 ;
      RECT 8.0200 0.8600 8.1300 0.9650 ;
      RECT 8.0200 0.9650 8.1100 1.6650 ;
  END
END POSTICG_X13B_A12TH

MACRO POSTICG_X16B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 10.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7300 ;
        RECT 0.6000 0.3200 0.6900 0.6150 ;
        RECT 1.1200 0.3200 1.2100 0.6150 ;
        RECT 1.6400 0.3200 1.7300 0.6150 ;
        RECT 2.1600 0.3200 2.2500 0.6150 ;
        RECT 2.6800 0.3200 2.7700 0.6500 ;
        RECT 5.0100 0.3200 5.1000 0.6600 ;
        RECT 5.5300 0.3200 5.6200 0.6600 ;
        RECT 6.0500 0.3200 6.1400 0.6600 ;
        RECT 6.5700 0.3200 6.6600 0.6750 ;
        RECT 7.0800 0.3200 7.1700 0.7300 ;
        RECT 8.0600 0.3200 8.1500 0.5350 ;
        RECT 9.8500 0.3200 9.9400 0.6650 ;
        RECT 10.3750 0.3200 10.4650 0.8850 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7900 1.2600 6.5550 1.3500 ;
        RECT 6.4550 1.3500 6.5550 1.8300 ;
        RECT 4.7900 1.2500 6.0650 1.2600 ;
        RECT 6.4550 1.8300 9.7400 1.9200 ;
        RECT 8.2350 1.1250 8.3250 1.8300 ;
        RECT 9.6500 1.1000 9.7400 1.8300 ;
    END
    ANTENNAGATEAREA 0.6012 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.0100 1.0400 10.4000 1.1500 ;
    END
    ANTENNAGATEAREA 0.1194 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9300 1.2400 7.4250 1.3600 ;
    END
    ANTENNAGATEAREA 0.144 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5900 0.9600 0.8100 1.3100 ;
        RECT 0.3400 1.3100 4.0700 1.5250 ;
        RECT 0.3400 0.7450 2.5100 0.9600 ;
        RECT 0.3400 1.5250 0.4300 1.7250 ;
        RECT 0.8600 1.5250 0.9500 1.7250 ;
        RECT 1.3800 1.5250 1.4700 1.7250 ;
        RECT 1.9000 1.5250 1.9900 1.7250 ;
        RECT 2.4200 1.5250 2.5100 1.7250 ;
        RECT 2.9400 1.5250 3.0300 1.7250 ;
        RECT 3.4600 1.5250 3.5500 1.7250 ;
        RECT 3.9800 1.5250 4.0700 1.7250 ;
        RECT 0.3400 0.5300 0.4300 0.7450 ;
        RECT 0.8600 0.5300 0.9500 0.7450 ;
        RECT 1.3800 0.5300 1.4700 0.7450 ;
        RECT 1.9000 0.5300 1.9900 0.7450 ;
        RECT 2.4200 0.4100 2.5100 0.7450 ;
    END
    ANTENNADIFFAREA 2.216 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 10.6450 2.7200 ;
        RECT 7.2700 2.0100 7.3600 2.0800 ;
        RECT 7.7900 2.0100 8.0800 2.0800 ;
        RECT 9.8500 1.7900 9.9400 2.0800 ;
        RECT 4.3450 1.7750 4.4350 2.0800 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
        RECT 1.1200 1.7700 1.2100 2.0800 ;
        RECT 1.6400 1.7700 1.7300 2.0800 ;
        RECT 2.1600 1.7700 2.2500 2.0800 ;
        RECT 2.6800 1.7700 2.7700 2.0800 ;
        RECT 3.2000 1.7700 3.2900 2.0800 ;
        RECT 3.7200 1.7700 3.8100 2.0800 ;
        RECT 4.9750 1.6400 5.0650 2.0800 ;
        RECT 5.4950 1.6400 5.5850 2.0800 ;
        RECT 6.0150 1.6400 6.1050 2.0800 ;
        RECT 10.3700 1.5700 10.4600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.4550 1.4600 6.3650 1.5500 ;
      RECT 6.2750 1.5500 6.3650 1.9000 ;
      RECT 2.9300 0.4100 3.0200 1.0650 ;
      RECT 3.4500 0.6600 3.5400 1.0650 ;
      RECT 3.9700 0.6600 4.0600 1.0650 ;
      RECT 4.7150 1.5500 4.8050 1.9150 ;
      RECT 4.4550 1.2000 4.5450 1.4600 ;
      RECT 1.5000 1.1100 4.5800 1.2000 ;
      RECT 2.9300 1.0650 4.5800 1.1100 ;
      RECT 4.4900 0.6600 4.5800 1.0650 ;
      RECT 5.2350 1.5500 5.3250 1.9000 ;
      RECT 5.7550 1.5500 5.8450 1.9000 ;
      RECT 4.7500 0.7700 6.4000 0.8600 ;
      RECT 5.7900 0.7500 6.4000 0.7700 ;
      RECT 6.3100 0.4100 6.4000 0.7500 ;
      RECT 4.7500 0.5700 4.8400 0.7700 ;
      RECT 3.1500 0.4800 4.8400 0.5700 ;
      RECT 3.1500 0.5700 3.3200 0.8100 ;
      RECT 3.6700 0.5700 3.8400 0.8100 ;
      RECT 4.1900 0.5700 4.3600 0.8100 ;
      RECT 5.2700 0.4100 5.3600 0.7700 ;
      RECT 5.7900 0.4100 5.8800 0.7500 ;
      RECT 6.8200 0.8200 7.4300 0.9100 ;
      RECT 7.3400 0.5700 7.4300 0.8200 ;
      RECT 7.3400 0.4800 7.9500 0.5700 ;
      RECT 7.8600 0.5700 7.9500 0.8350 ;
      RECT 6.8200 0.4800 6.9100 0.8200 ;
      RECT 6.6650 1.6500 8.0950 1.7400 ;
      RECT 8.0050 1.3750 8.0950 1.6500 ;
      RECT 7.6000 0.7600 7.6900 1.6500 ;
      RECT 6.6650 1.0750 6.7550 1.6500 ;
      RECT 5.0850 0.9850 6.7550 1.0750 ;
      RECT 8.5600 1.6500 9.2100 1.7400 ;
      RECT 8.6050 1.0350 8.6950 1.6500 ;
      RECT 9.1200 0.7550 9.2100 1.6500 ;
      RECT 7.7850 0.9450 8.6950 1.0350 ;
      RECT 9.0650 0.6600 9.2750 0.7550 ;
      RECT 8.6050 0.4100 8.6950 0.9450 ;
      RECT 7.7850 1.0350 7.8750 1.3000 ;
      RECT 9.4500 1.1300 9.5400 1.6300 ;
      RECT 9.4200 0.9200 9.5400 1.1300 ;
      RECT 9.4500 0.6800 9.5400 0.9200 ;
      RECT 10.1100 1.5900 10.2000 1.9300 ;
      RECT 9.8300 1.5000 10.2000 1.5900 ;
      RECT 9.6700 0.8100 10.2050 0.9000 ;
      RECT 10.1150 0.4400 10.2050 0.8100 ;
      RECT 9.8300 0.9000 9.9200 1.5000 ;
      RECT 9.6700 0.5700 9.7600 0.8100 ;
      RECT 8.8650 0.4800 9.7600 0.5700 ;
      RECT 8.8650 0.5700 8.9550 1.4250 ;
      RECT 8.8650 0.4250 8.9550 0.4800 ;
      RECT 8.8200 1.4250 8.9900 1.5150 ;
  END
END POSTICG_X16B_A12TH

MACRO POSTICG_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.7000 ;
        RECT 1.4900 0.3200 1.7000 0.7200 ;
        RECT 2.6300 0.3200 2.8400 0.3900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0350 2.9550 1.3750 ;
        RECT 2.6550 1.3750 2.9550 1.4650 ;
        RECT 2.6550 1.4650 2.7450 1.8300 ;
        RECT 0.8500 1.8300 2.7450 1.9200 ;
        RECT 2.2750 1.3500 2.3650 1.8300 ;
        RECT 0.8500 1.3400 0.9400 1.8300 ;
        RECT 1.8650 1.2600 2.3650 1.3500 ;
        RECT 0.7900 1.1700 0.9400 1.3400 ;
        RECT 1.8650 1.1100 1.9550 1.2600 ;
    END
    ANTENNAGATEAREA 0.0804 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6350 0.8300 2.7500 1.2050 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END E

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0100 1.5500 1.1750 ;
        RECT 1.2300 1.1750 1.5500 1.2650 ;
    END
    ANTENNAGATEAREA 0.0258 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7800 0.1500 1.2900 ;
        RECT 0.0500 1.2900 0.1750 1.7200 ;
        RECT 0.0500 0.6350 0.1750 0.7800 ;
        RECT 0.0750 0.4100 0.1750 0.6350 ;
    END
    ANTENNADIFFAREA 0.2184 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.4500 2.0100 1.6200 2.0800 ;
        RECT 2.8300 1.9550 2.9200 2.0800 ;
        RECT 0.2800 1.6550 0.4900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3100 0.7900 0.9050 0.8800 ;
      RECT 0.8150 0.5600 0.9050 0.7900 ;
      RECT 0.6500 1.5350 0.7400 1.8050 ;
      RECT 0.3100 1.4450 0.7400 1.5350 ;
      RECT 0.3100 1.1400 0.4000 1.4450 ;
      RECT 0.2400 0.9300 0.4000 1.1400 ;
      RECT 0.3100 0.8800 0.4000 0.9300 ;
      RECT 1.0300 1.6300 1.5950 1.7200 ;
      RECT 1.5050 1.3750 1.5950 1.6300 ;
      RECT 1.0300 1.0600 1.1200 1.6300 ;
      RECT 0.5150 0.9700 1.1200 1.0600 ;
      RECT 1.0300 0.7150 1.1200 0.9700 ;
      RECT 1.0300 0.6250 1.2350 0.7150 ;
      RECT 0.5150 1.0600 0.6050 1.3500 ;
      RECT 1.9750 1.6400 2.1650 1.7200 ;
      RECT 1.6850 1.6300 2.1650 1.6400 ;
      RECT 1.6850 1.5500 2.0650 1.6300 ;
      RECT 1.2100 0.8300 2.0400 0.9200 ;
      RECT 1.9500 0.7500 2.0400 0.8300 ;
      RECT 1.9500 0.6600 2.1700 0.7500 ;
      RECT 1.6850 0.9200 1.7750 1.5500 ;
      RECT 1.2100 0.9200 1.3000 1.0550 ;
      RECT 2.4550 0.7500 2.5450 1.7100 ;
      RECT 2.2900 0.6600 2.5450 0.7500 ;
      RECT 3.0300 1.5550 3.1550 1.7650 ;
      RECT 3.0650 0.7750 3.1550 1.5550 ;
      RECT 3.0300 0.5700 3.1550 0.7750 ;
      RECT 2.0750 0.4800 3.1550 0.5700 ;
      RECT 2.0750 0.4100 2.2850 0.4800 ;
  END
END POSTICG_X1B_A12TH

MACRO POSTICG_X1P2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.4900 0.3200 0.5800 0.8200 ;
        RECT 1.6950 0.3200 1.7850 0.6850 ;
        RECT 3.0300 0.3200 3.2400 0.3900 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.6200 ;
        RECT 0.0500 1.6200 0.4400 1.7200 ;
        RECT 0.0500 0.8500 0.3250 0.9500 ;
        RECT 0.3400 1.7200 0.4400 1.9900 ;
        RECT 0.2250 0.4100 0.3250 0.8500 ;
    END
    ANTENNADIFFAREA 0.198 ;
  END ECK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0400 0.8100 3.1500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.6550 2.9500 1.8300 ;
        RECT 1.1800 1.8300 2.9500 1.9200 ;
        RECT 2.8500 1.5650 3.1300 1.6550 ;
        RECT 1.1800 1.5100 1.2700 1.8300 ;
        RECT 2.4500 1.2550 2.5400 1.8300 ;
        RECT 3.0400 1.4950 3.1300 1.5650 ;
        RECT 1.0600 1.4200 1.2700 1.5100 ;
        RECT 2.2200 1.1650 2.7700 1.2550 ;
        RECT 3.0400 1.4050 3.3600 1.4950 ;
        RECT 2.2200 0.9550 2.3100 1.1650 ;
        RECT 3.2700 1.2850 3.3600 1.4050 ;
    END
    ANTENNAGATEAREA 0.0867 ;
  END CK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5700 1.0500 1.8950 1.1500 ;
        RECT 1.5700 0.9550 1.6700 1.0500 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END SEN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.0450 1.8400 0.2150 2.0800 ;
        RECT 0.6050 1.7500 0.6950 2.0800 ;
        RECT 3.0400 1.7450 3.2500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.9150 1.6900 1.0050 1.9600 ;
      RECT 0.8600 1.6000 1.0050 1.6900 ;
      RECT 0.8600 1.5000 0.9500 1.6000 ;
      RECT 0.2400 1.4100 0.9500 1.5000 ;
      RECT 0.5350 1.0000 0.6250 1.4100 ;
      RECT 0.5350 0.9100 1.0400 1.0000 ;
      RECT 0.9500 0.4400 1.0400 0.9100 ;
      RECT 1.1300 1.2400 1.9300 1.3300 ;
      RECT 1.8350 1.3300 1.9300 1.4550 ;
      RECT 1.4750 1.3300 1.5650 1.7400 ;
      RECT 1.1300 1.1900 1.2200 1.2400 ;
      RECT 0.7350 1.1000 1.2200 1.1900 ;
      RECT 1.1300 0.6450 1.2200 1.1000 ;
      RECT 1.1300 0.5550 1.3550 0.6450 ;
      RECT 0.7350 1.1900 0.8250 1.2900 ;
      RECT 2.2500 1.6400 2.3400 1.7400 ;
      RECT 2.0200 1.5500 2.3400 1.6400 ;
      RECT 1.3200 0.7750 2.4200 0.8650 ;
      RECT 2.3300 0.5650 2.4200 0.7750 ;
      RECT 2.0200 0.8650 2.1100 1.5500 ;
      RECT 1.3200 0.8650 1.4100 0.9600 ;
      RECT 2.6500 1.3850 2.9500 1.4750 ;
      RECT 2.8600 0.7500 2.9500 1.3850 ;
      RECT 2.7100 0.6600 2.9500 0.7500 ;
      RECT 2.6500 1.4750 2.7400 1.7400 ;
      RECT 3.4250 1.5850 3.5400 1.7950 ;
      RECT 3.4500 0.7950 3.5400 1.5850 ;
      RECT 3.4250 0.5700 3.5400 0.7950 ;
      RECT 2.5100 0.4800 3.5400 0.5700 ;
      RECT 2.5100 0.5700 2.6000 1.0250 ;
  END
END POSTICG_X1P2B_A12TH

MACRO POSTICG_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.7650 ;
        RECT 1.6500 0.3200 1.8600 0.6250 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4500 0.4350 1.5500 ;
        RECT 0.3350 1.5500 0.4350 1.9750 ;
        RECT 0.0500 0.9800 0.1500 1.4500 ;
        RECT 0.0500 0.9000 0.1750 0.9800 ;
        RECT 0.0750 0.5400 0.1750 0.9000 ;
    END
    ANTENNADIFFAREA 0.2286 ;
  END ECK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9550 1.0350 3.3200 1.1550 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0000 1.4600 2.1500 1.5500 ;
        RECT 2.0500 1.5500 2.1500 1.8300 ;
        RECT 1.0000 1.3850 1.1950 1.4600 ;
        RECT 2.0500 1.8300 3.0450 1.9200 ;
        RECT 2.9550 1.4800 3.0450 1.8300 ;
        RECT 2.5950 1.1900 2.6850 1.8300 ;
        RECT 2.9550 1.3800 3.3400 1.4800 ;
        RECT 2.2650 1.1000 2.6850 1.1900 ;
        RECT 3.2500 1.3000 3.3400 1.3800 ;
        RECT 2.2650 0.8500 2.3550 1.1000 ;
    END
    ANTENNAGATEAREA 0.0933 ;
  END CK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 1.0500 1.7050 1.1500 ;
        RECT 1.5350 0.9000 1.7050 1.0500 ;
    END
    ANTENNAGATEAREA 0.0294 ;
  END SEN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.6000 2.0000 0.6900 2.0800 ;
        RECT 1.2100 1.8200 1.3800 2.0800 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 1.8500 1.6650 1.9400 2.0800 ;
        RECT 3.1350 1.5900 3.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5450 1.0700 0.6350 1.1500 ;
      RECT 0.5450 1.3600 0.6350 1.8200 ;
      RECT 0.5450 0.9800 1.0500 1.0700 ;
      RECT 0.5450 1.8200 1.0700 1.9100 ;
      RECT 0.9600 0.5400 1.0500 0.9800 ;
      RECT 0.9800 1.9100 1.0700 1.9900 ;
      RECT 0.3650 1.1500 0.6350 1.3600 ;
      RECT 1.1900 0.7150 1.9350 0.8050 ;
      RECT 1.8450 0.8050 1.9350 0.9850 ;
      RECT 1.5900 1.7300 1.6800 1.8900 ;
      RECT 0.8000 1.6400 1.6800 1.7300 ;
      RECT 0.8000 1.4600 0.8900 1.6400 ;
      RECT 0.7300 1.2500 0.8900 1.4600 ;
      RECT 0.8000 1.1600 1.2800 1.2500 ;
      RECT 1.1900 0.8050 1.2800 1.1600 ;
      RECT 1.1900 0.5150 1.2800 0.7150 ;
      RECT 2.2950 1.6450 2.4850 1.7350 ;
      RECT 2.2950 1.3700 2.3850 1.6450 ;
      RECT 1.4250 1.2800 2.3850 1.3700 ;
      RECT 2.0250 0.6500 2.3900 0.7400 ;
      RECT 2.3000 0.5450 2.3900 0.6500 ;
      RECT 2.0250 0.7400 2.1150 1.2800 ;
      RECT 2.7750 0.7600 2.8650 1.7200 ;
      RECT 2.6950 0.6700 2.8650 0.7600 ;
      RECT 3.4300 1.5650 3.5300 1.7750 ;
      RECT 3.4400 0.9000 3.5300 1.5650 ;
      RECT 2.9550 0.8100 3.5300 0.9000 ;
      RECT 3.4300 0.5950 3.5300 0.8100 ;
      RECT 2.4950 0.5800 2.5850 0.9000 ;
      RECT 2.4950 0.5600 2.7900 0.5800 ;
      RECT 2.4950 0.9000 2.6850 0.9900 ;
      RECT 2.9550 0.5600 3.0450 0.8100 ;
      RECT 2.4950 0.4900 3.0450 0.5600 ;
      RECT 2.6950 0.4700 3.0450 0.4900 ;
  END
END POSTICG_X1P4B_A12TH

MACRO POSTICG_X1P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 1.5950 0.3200 1.8050 0.5750 ;
        RECT 3.0950 0.3200 3.1850 0.7000 ;
    END
  END VSS

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3000 0.8500 1.6400 0.9500 ;
        RECT 1.5400 0.9500 1.6400 1.1200 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4500 0.4050 1.5500 ;
        RECT 0.3150 1.5500 0.4050 1.6000 ;
        RECT 0.0500 0.9900 0.1500 1.4500 ;
        RECT 0.3150 1.6000 0.4350 1.6900 ;
        RECT 0.0500 0.8650 0.1750 0.9900 ;
        RECT 0.3350 1.6900 0.4350 1.9700 ;
        RECT 0.0750 0.5400 0.1750 0.8650 ;
    END
    ANTENNADIFFAREA 0.2772 ;
  END ECK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9200 1.0450 3.3200 1.1550 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8700 1.1500 1.3900 ;
        RECT 1.0500 1.3900 1.9100 1.4800 ;
        RECT 1.8200 1.4800 2.1800 1.5700 ;
        RECT 2.0900 1.5700 2.1800 1.8300 ;
        RECT 2.0900 1.8300 3.0800 1.9200 ;
        RECT 2.9900 1.5150 3.0800 1.8300 ;
        RECT 2.5500 1.1950 2.6400 1.8300 ;
        RECT 2.9900 1.4150 3.3400 1.5150 ;
        RECT 2.2200 1.1050 2.6400 1.1950 ;
        RECT 3.2500 1.3050 3.3400 1.4150 ;
        RECT 2.2200 0.9300 2.3100 1.1050 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.6000 2.0000 0.6900 2.0800 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 1.2600 1.7500 1.3600 2.0800 ;
        RECT 1.7850 1.6600 1.9950 2.0800 ;
        RECT 3.1700 1.6250 3.2600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6050 1.7500 1.1300 1.8400 ;
      RECT 0.6050 1.5100 0.6950 1.7500 ;
      RECT 0.4950 1.4200 0.6950 1.5100 ;
      RECT 0.4950 1.2950 0.5850 1.4200 ;
      RECT 0.2500 1.2050 0.5850 1.2950 ;
      RECT 0.4950 0.5700 0.5850 1.2050 ;
      RECT 0.4950 0.4800 1.0050 0.5700 ;
      RECT 0.8050 0.6700 1.9300 0.7600 ;
      RECT 1.8400 0.7600 1.9300 0.9500 ;
      RECT 1.5850 1.6600 1.6750 1.8500 ;
      RECT 0.8050 1.5700 1.6750 1.6600 ;
      RECT 0.8050 1.2800 0.8950 1.5700 ;
      RECT 0.7350 1.0700 0.8950 1.2800 ;
      RECT 0.8050 0.7600 0.8950 1.0700 ;
      RECT 1.1600 0.4900 1.2500 0.6700 ;
      RECT 2.2700 1.6300 2.4600 1.7200 ;
      RECT 2.2700 1.3900 2.3600 1.6300 ;
      RECT 2.0400 1.3000 2.3600 1.3900 ;
      RECT 2.0400 0.7200 2.3400 0.8100 ;
      RECT 2.2500 0.5200 2.3400 0.7200 ;
      RECT 1.4400 1.2100 2.1300 1.3000 ;
      RECT 2.0400 0.8100 2.1300 1.2100 ;
      RECT 2.7300 1.6300 2.9000 1.7200 ;
      RECT 2.7300 0.7500 2.8200 1.6300 ;
      RECT 2.6500 0.6600 2.8200 0.7500 ;
      RECT 3.4300 1.5700 3.5300 1.8150 ;
      RECT 3.4400 0.9000 3.5300 1.5700 ;
      RECT 2.9150 0.8100 3.5300 0.9000 ;
      RECT 3.4300 0.5850 3.5300 0.8100 ;
      RECT 2.4500 0.5700 2.5400 0.9050 ;
      RECT 2.4500 0.9050 2.6400 0.9950 ;
      RECT 2.9150 0.5700 3.0050 0.8100 ;
      RECT 2.4500 0.4800 3.0050 0.5700 ;
  END
END POSTICG_X1P7B_A12TH

MACRO POSTICG_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7500 ;
        RECT 0.6000 0.3200 0.6900 0.7500 ;
        RECT 1.7100 0.3200 1.9200 0.5200 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2500 0.4300 1.3500 ;
        RECT 0.3400 1.3500 0.4300 1.7200 ;
        RECT 0.0500 0.9500 0.1500 1.2500 ;
        RECT 0.0500 0.8500 0.4300 0.9500 ;
        RECT 0.3400 0.4100 0.4300 0.8500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6450 0.8100 1.7850 1.1350 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9550 1.0400 3.3150 1.1600 ;
    END
    ANTENNAGATEAREA 0.033 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.2500 1.1950 1.4200 ;
        RECT 1.0100 1.4200 2.1500 1.5100 ;
        RECT 2.0500 1.5100 2.1500 1.8300 ;
        RECT 2.0500 1.8300 3.0800 1.9200 ;
        RECT 2.9900 1.5150 3.0800 1.8300 ;
        RECT 2.5500 1.1500 2.6400 1.8300 ;
        RECT 2.9900 1.4250 3.3400 1.5150 ;
        RECT 2.2550 1.0600 2.6400 1.1500 ;
        RECT 3.2500 1.3050 3.3400 1.4250 ;
        RECT 2.2550 0.9100 2.3450 1.0600 ;
    END
    ANTENNAGATEAREA 0.1137 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.6000 2.0200 0.6900 2.0800 ;
        RECT 1.2500 1.7800 1.3400 2.0800 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 3.1700 1.6250 3.2600 2.0800 ;
        RECT 1.8650 1.6200 1.9550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5350 1.8100 1.1400 1.9000 ;
      RECT 0.5350 0.8900 1.1500 0.9800 ;
      RECT 1.0600 0.4750 1.1500 0.8900 ;
      RECT 0.5350 1.1500 0.6250 1.8100 ;
      RECT 0.3000 1.0600 0.6250 1.1500 ;
      RECT 0.5350 0.9800 0.6250 1.0600 ;
      RECT 1.2400 0.6100 1.9650 0.7000 ;
      RECT 1.8750 0.7000 1.9650 0.9150 ;
      RECT 0.7650 1.1600 0.8550 1.6000 ;
      RECT 1.6000 1.6900 1.6900 1.8650 ;
      RECT 0.7650 1.6000 1.6900 1.6900 ;
      RECT 0.7650 1.0700 1.3300 1.1600 ;
      RECT 1.2400 0.7000 1.3300 1.0700 ;
      RECT 1.2400 0.5700 1.4000 0.6100 ;
      RECT 1.3100 0.4500 1.4000 0.5700 ;
      RECT 2.2700 1.6300 2.4600 1.7200 ;
      RECT 2.2700 1.3300 2.3600 1.6300 ;
      RECT 1.4350 1.2400 2.3600 1.3300 ;
      RECT 2.0550 0.6100 2.3850 0.7000 ;
      RECT 2.2950 0.4950 2.3850 0.6100 ;
      RECT 2.0550 0.7000 2.1450 1.2400 ;
      RECT 2.7300 1.6300 2.9000 1.7200 ;
      RECT 2.7550 0.7500 2.8450 1.6300 ;
      RECT 2.6750 0.6600 2.8450 0.7500 ;
      RECT 3.4300 1.5850 3.5300 1.8150 ;
      RECT 3.4400 0.7950 3.5300 1.5850 ;
      RECT 3.4300 0.5700 3.5300 0.7950 ;
      RECT 2.4750 0.4800 3.5300 0.5700 ;
      RECT 2.4750 0.5700 2.5650 0.8800 ;
      RECT 2.4750 0.8800 2.6450 0.9700 ;
  END
END POSTICG_X2B_A12TH

MACRO POSTICG_X2P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.2000 0.3200 0.2900 0.6800 ;
        RECT 0.7500 0.3200 0.8500 0.4500 ;
        RECT 1.8950 0.3200 2.1050 0.4850 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 0.6950 1.5500 ;
        RECT 0.0750 1.5500 0.1750 1.8700 ;
        RECT 0.5950 1.5500 0.6950 1.8700 ;
        RECT 0.0750 0.9500 0.1750 1.4500 ;
        RECT 0.0750 0.8500 0.5550 0.9500 ;
        RECT 0.4550 0.4100 0.5550 0.8500 ;
    END
    ANTENNADIFFAREA 0.3876 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.8100 1.9900 0.9500 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1550 1.0350 3.5250 1.1550 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END E

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.3400 1.8400 0.4300 2.0800 ;
        RECT 1.4950 1.7700 1.5850 2.0800 ;
        RECT 2.0400 1.6100 2.2500 2.0800 ;
        RECT 3.3350 1.5300 3.4250 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.0500 1.3900 1.2500 ;
        RECT 1.2100 1.2500 2.1850 1.3500 ;
        RECT 2.0950 1.3500 2.1850 1.4300 ;
        RECT 2.0950 1.4300 2.4850 1.5200 ;
        RECT 2.3950 1.5200 2.4850 1.8300 ;
        RECT 2.3950 1.8300 3.2250 1.9200 ;
        RECT 3.1350 1.4400 3.2250 1.8300 ;
        RECT 2.7750 1.1600 2.8650 1.8300 ;
        RECT 3.1350 1.3500 3.5400 1.4400 ;
        RECT 2.4750 1.0700 2.8650 1.1600 ;
        RECT 3.4500 1.2600 3.5400 1.3500 ;
        RECT 2.4750 0.8150 2.5650 1.0700 ;
    END
    ANTENNAGATEAREA 0.1299 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 1.2350 1.7100 1.3250 1.9900 ;
      RECT 0.8000 1.6200 1.3250 1.7100 ;
      RECT 0.8000 0.6900 1.3100 0.7800 ;
      RECT 1.2200 0.4100 1.3100 0.6900 ;
      RECT 0.8000 1.3300 0.8900 1.6200 ;
      RECT 0.4150 1.2400 0.8900 1.3300 ;
      RECT 0.8000 0.7800 0.8900 1.2400 ;
      RECT 1.4300 0.6100 2.1850 0.7000 ;
      RECT 2.0950 0.7000 2.1850 0.9550 ;
      RECT 1.8400 1.5300 1.9300 1.7750 ;
      RECT 0.9800 1.4400 1.9300 1.5300 ;
      RECT 0.9800 0.9600 1.0700 1.4400 ;
      RECT 0.9800 0.8700 1.5200 0.9600 ;
      RECT 1.4300 0.7000 1.5200 0.8700 ;
      RECT 1.4300 0.5400 1.5600 0.6100 ;
      RECT 1.4700 0.4200 1.5600 0.5400 ;
      RECT 2.5950 1.3400 2.6850 1.7200 ;
      RECT 2.2750 1.2500 2.6850 1.3400 ;
      RECT 2.2750 0.6100 2.5850 0.7000 ;
      RECT 2.4950 0.4850 2.5850 0.6100 ;
      RECT 2.2750 1.1600 2.3650 1.2500 ;
      RECT 1.5950 1.0700 2.3650 1.1600 ;
      RECT 2.2750 0.7000 2.3650 1.0700 ;
      RECT 2.9550 0.7500 3.0450 1.7200 ;
      RECT 2.8750 0.6600 3.0450 0.7500 ;
      RECT 3.6300 1.5400 3.7500 1.7450 ;
      RECT 3.6600 0.7750 3.7500 1.5400 ;
      RECT 3.6300 0.5700 3.7500 0.7750 ;
      RECT 2.6750 0.4800 3.7500 0.5700 ;
      RECT 2.6750 0.5700 2.7650 0.8900 ;
      RECT 2.6750 0.8900 2.8450 0.9800 ;
  END
END POSTICG_X2P5B_A12TH

MACRO POSTICG_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.5600 0.3200 0.6500 0.7400 ;
        RECT 1.2750 0.3200 1.6450 0.4500 ;
        RECT 2.4750 0.3200 2.5650 0.7000 ;
        RECT 3.9500 0.3200 4.0400 0.6950 ;
    END
  END VSS

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.5650 1.4450 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SEN

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9900 1.2500 1.6100 1.3500 ;
        RECT 0.9900 1.3500 1.0900 1.6350 ;
        RECT 1.5200 1.3500 1.6100 1.6600 ;
        RECT 0.9900 0.7600 1.0900 1.2500 ;
    END
    ANTENNADIFFAREA 0.51815 ;
  END ECK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7700 1.0400 4.1250 1.1600 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7700 1.4900 4.1650 1.5900 ;
        RECT 3.7700 1.5900 3.8600 1.8300 ;
        RECT 4.0500 1.4100 4.1650 1.4900 ;
        RECT 2.9300 1.8300 3.8600 1.9200 ;
        RECT 3.3700 1.2250 3.4600 1.8300 ;
        RECT 2.9300 1.1500 3.0200 1.8300 ;
        RECT 2.5200 1.1300 3.0200 1.1500 ;
        RECT 2.5200 1.1500 2.6100 1.2350 ;
        RECT 1.9550 1.0300 3.0200 1.1300 ;
    END
    ANTENNAGATEAREA 0.1467 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 1.2600 1.9500 1.3500 2.0800 ;
        RECT 0.0800 1.7150 0.1700 2.0800 ;
        RECT 0.6000 1.7150 0.6900 2.0800 ;
        RECT 3.9700 1.6800 4.0600 2.0800 ;
        RECT 2.0300 1.4850 2.1200 2.0800 ;
        RECT 2.6250 1.4850 2.7150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8000 1.7500 1.8600 1.8400 ;
      RECT 0.3400 1.6250 0.4300 1.9500 ;
      RECT 0.0450 0.7400 0.1350 1.5350 ;
      RECT 0.0450 0.6050 0.2250 0.7400 ;
      RECT 0.0550 0.4300 0.2250 0.6050 ;
      RECT 0.8000 1.6250 0.8900 1.7500 ;
      RECT 0.0450 1.5350 0.8900 1.6250 ;
      RECT 2.3650 1.3950 2.4550 1.7900 ;
      RECT 1.7300 1.3050 2.4550 1.3950 ;
      RECT 1.7300 0.7500 2.0450 0.8400 ;
      RECT 1.9550 0.6600 2.1550 0.7500 ;
      RECT 1.7300 1.1600 1.8200 1.3050 ;
      RECT 1.2000 1.0700 1.8200 1.1600 ;
      RECT 1.7300 0.8400 1.8200 1.0700 ;
      RECT 3.1900 1.5600 3.2800 1.6950 ;
      RECT 3.1100 1.4700 3.2800 1.5600 ;
      RECT 3.1100 0.9000 3.2000 1.4700 ;
      RECT 2.2750 0.8100 3.2000 0.9000 ;
      RECT 3.1100 0.5050 3.2000 0.8100 ;
      RECT 0.2250 0.9400 0.3150 1.2400 ;
      RECT 0.7500 0.5700 1.8650 0.6500 ;
      RECT 0.7500 0.6500 0.8400 0.8500 ;
      RECT 0.2250 0.8500 0.8400 0.9400 ;
      RECT 2.2750 0.5700 2.3650 0.8100 ;
      RECT 0.7500 0.5600 2.3650 0.5700 ;
      RECT 1.7750 0.4800 2.3650 0.5600 ;
      RECT 3.5700 0.7700 3.6600 1.7400 ;
      RECT 3.4900 0.6800 3.6600 0.7700 ;
      RECT 4.2300 1.7700 4.3200 1.8900 ;
      RECT 4.2300 1.6800 4.3450 1.7700 ;
      RECT 4.2550 0.9000 4.3450 1.6800 ;
      RECT 3.7500 0.8100 4.3450 0.9000 ;
      RECT 4.2300 0.6250 4.3450 0.8100 ;
      RECT 4.2300 0.5050 4.3200 0.6250 ;
      RECT 3.2900 0.5700 3.3800 1.0950 ;
      RECT 3.7500 0.5700 3.8400 0.8100 ;
      RECT 3.2900 0.4800 3.8400 0.5700 ;
  END
END POSTICG_X3B_A12TH

MACRO POSTICG_X3P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.6650 ;
        RECT 0.9250 0.3200 1.0150 0.4850 ;
        RECT 1.9400 0.3200 2.0300 0.6000 ;
        RECT 2.5950 0.3200 2.7850 0.6050 ;
        RECT 3.9350 0.3200 4.0250 0.6650 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.4500 0.9500 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8200 ;
        RECT 0.8600 1.5500 0.9500 1.8200 ;
        RECT 0.1000 0.9500 0.2000 1.4500 ;
        RECT 0.1000 0.8500 0.7150 0.9500 ;
        RECT 0.6250 0.4250 0.7150 0.8500 ;
        RECT 0.1000 0.4100 0.1950 0.8500 ;
    END
    ANTENNADIFFAREA 0.57 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8600 1.0200 2.2550 1.1500 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7550 1.0350 4.1150 1.1600 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 1.0350 1.7500 1.1500 ;
        RECT 1.6500 1.1500 1.7500 1.2600 ;
        RECT 1.6500 1.2600 2.2400 1.3500 ;
        RECT 2.1500 1.3500 2.2400 1.4700 ;
        RECT 2.1500 1.4700 2.9500 1.5700 ;
        RECT 2.8500 1.5700 2.9500 1.8300 ;
        RECT 2.8500 1.8300 3.8800 1.9200 ;
        RECT 3.7900 1.4850 3.8800 1.8300 ;
        RECT 3.3500 1.1800 3.4400 1.8300 ;
        RECT 3.7900 1.3850 4.1650 1.4850 ;
        RECT 3.0200 1.0900 3.4400 1.1800 ;
        RECT 4.0750 1.3000 4.1650 1.3850 ;
        RECT 3.0200 0.9400 3.1100 1.0900 ;
    END
    ANTENNAGATEAREA 0.1563 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 1.1300 2.0200 1.2200 2.0800 ;
        RECT 0.0800 1.7650 0.1700 2.0800 ;
        RECT 0.6000 1.7650 0.6900 2.0800 ;
        RECT 1.7800 1.7500 1.8700 2.0800 ;
        RECT 2.4900 1.7500 2.5800 2.0800 ;
        RECT 3.9700 1.5950 4.0600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.5000 1.7100 1.5900 1.9900 ;
      RECT 1.0400 1.6200 1.5900 1.7100 ;
      RECT 0.9650 0.6100 1.5700 0.7000 ;
      RECT 1.4800 0.4650 1.5700 0.6100 ;
      RECT 1.0400 1.2750 1.1300 1.6200 ;
      RECT 0.4700 1.1850 1.1300 1.2750 ;
      RECT 0.9650 0.7000 1.0550 1.1850 ;
      RECT 1.1450 0.8150 2.7300 0.9050 ;
      RECT 1.2200 1.0300 1.3100 1.4400 ;
      RECT 1.1450 0.9050 1.3100 1.0300 ;
      RECT 2.4000 0.4300 2.4900 0.8150 ;
      RECT 2.1750 1.7500 2.2650 1.9900 ;
      RECT 1.9700 1.6600 2.2650 1.7500 ;
      RECT 1.9700 1.5300 2.0600 1.6600 ;
      RECT 1.2200 1.4400 2.0600 1.5300 ;
      RECT 3.0700 1.6300 3.2600 1.7200 ;
      RECT 3.0700 1.3600 3.1600 1.6300 ;
      RECT 2.3300 1.2700 3.1600 1.3600 ;
      RECT 2.8200 0.7400 3.1850 0.8300 ;
      RECT 3.0950 0.4550 3.1850 0.7400 ;
      RECT 2.8200 0.8300 2.9100 1.2700 ;
      RECT 3.5300 1.6250 3.7000 1.7150 ;
      RECT 3.5550 0.7500 3.6450 1.6250 ;
      RECT 3.4750 0.6600 3.6450 0.7500 ;
      RECT 4.2300 1.6650 4.3200 1.8050 ;
      RECT 4.2300 1.5750 4.3450 1.6650 ;
      RECT 4.2550 0.8950 4.3450 1.5750 ;
      RECT 3.7350 0.8050 4.3450 0.8950 ;
      RECT 4.2300 0.7150 4.3450 0.8050 ;
      RECT 4.2300 0.4550 4.3200 0.7150 ;
      RECT 3.2750 0.5700 3.3650 0.8900 ;
      RECT 3.2750 0.8900 3.4650 0.9800 ;
      RECT 3.7350 0.5700 3.8250 0.8050 ;
      RECT 3.2750 0.4800 3.8250 0.5700 ;
  END
END POSTICG_X3P5B_A12TH

MACRO POSTICG_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.4400 0.3200 0.5300 0.6600 ;
        RECT 0.9950 0.3200 1.0850 0.5950 ;
        RECT 2.0450 0.3200 2.1350 0.5700 ;
        RECT 2.7550 0.3200 2.9250 0.5750 ;
        RECT 4.1500 0.3200 4.2400 0.6200 ;
    END
  END VSS

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 0.8500 2.5200 0.9500 ;
        RECT 2.2100 0.9500 2.3000 1.1600 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9600 1.0400 4.3300 1.1600 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5300 1.2500 2.8700 1.3500 ;
        RECT 2.7700 1.3500 2.8700 1.4450 ;
        RECT 1.5300 1.1850 1.9000 1.2500 ;
        RECT 2.7700 1.4450 3.2400 1.5350 ;
        RECT 3.1500 1.5350 3.2400 1.8300 ;
        RECT 3.1500 1.8300 4.0800 1.9200 ;
        RECT 3.9900 1.5350 4.0800 1.8300 ;
        RECT 3.5800 1.1750 3.6700 1.8300 ;
        RECT 3.9900 1.4350 4.3400 1.5350 ;
        RECT 3.1700 1.0850 3.6700 1.1750 ;
        RECT 4.2500 1.3000 4.3400 1.4350 ;
        RECT 3.1700 0.9650 3.2600 1.0850 ;
    END
    ANTENNAGATEAREA 0.1803 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 0.9500 1.3500 ;
        RECT 0.3350 1.3500 0.4350 1.7000 ;
        RECT 0.8500 1.3500 0.9500 1.7000 ;
        RECT 0.2500 0.9500 0.3500 1.2500 ;
        RECT 0.1750 0.8500 0.7950 0.9500 ;
        RECT 0.6950 0.4850 0.7950 0.8500 ;
        RECT 0.1750 0.4700 0.2750 0.8500 ;
    END
    ANTENNADIFFAREA 0.63 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 1.1200 2.0400 1.2100 2.0800 ;
        RECT 1.7550 1.8350 1.8450 2.0800 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
        RECT 4.1700 1.6450 4.2600 2.0800 ;
        RECT 2.2800 1.6350 2.3700 2.0800 ;
        RECT 2.8450 1.6300 2.9350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0400 1.6550 2.1050 1.7450 ;
      RECT 2.0150 1.7450 2.1050 1.8750 ;
      RECT 1.4950 1.7450 1.5850 1.8750 ;
      RECT 1.0400 0.7000 1.6500 0.7900 ;
      RECT 1.5600 0.4200 1.6500 0.7000 ;
      RECT 1.0400 1.1600 1.1300 1.6550 ;
      RECT 0.5000 1.0700 1.1300 1.1600 ;
      RECT 1.0400 0.7900 1.1300 1.0700 ;
      RECT 1.9450 0.6650 2.9000 0.7550 ;
      RECT 2.8100 0.7550 2.9000 0.8900 ;
      RECT 1.3250 1.0900 1.4150 1.4550 ;
      RECT 1.2200 1.0750 1.4150 1.0900 ;
      RECT 1.2200 0.9000 1.3100 0.9850 ;
      RECT 1.2200 0.9850 2.0350 1.0750 ;
      RECT 1.9450 0.7550 2.0350 0.9850 ;
      RECT 2.5400 1.5450 2.6300 1.9900 ;
      RECT 1.3250 1.4550 2.6300 1.5450 ;
      RECT 2.5450 0.4250 2.6350 0.6650 ;
      RECT 3.3800 1.3550 3.4700 1.7400 ;
      RECT 2.9900 1.2650 3.4700 1.3550 ;
      RECT 2.9900 0.7150 3.4000 0.8050 ;
      RECT 3.3100 0.4300 3.4000 0.7150 ;
      RECT 2.9900 1.1500 3.0800 1.2650 ;
      RECT 2.5500 1.0350 3.0800 1.1500 ;
      RECT 2.9900 0.8050 3.0800 1.0350 ;
      RECT 3.7800 0.7500 3.8700 1.7400 ;
      RECT 3.7000 0.6600 3.8700 0.7500 ;
      RECT 4.4300 1.6300 4.5300 1.8200 ;
      RECT 4.4400 0.8200 4.5300 1.6300 ;
      RECT 3.9700 0.7300 4.5300 0.8200 ;
      RECT 4.4300 0.4200 4.5300 0.7300 ;
      RECT 3.4900 0.5700 3.5800 0.8850 ;
      RECT 3.4900 0.8850 3.6800 0.9750 ;
      RECT 3.9700 0.5700 4.0600 0.7300 ;
      RECT 3.4900 0.4800 4.0600 0.5700 ;
  END
END POSTICG_X4B_A12TH

MACRO POSTICG_X5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.6550 0.3200 0.7450 0.6000 ;
        RECT 1.2250 0.3200 1.3150 0.6400 ;
        RECT 2.2750 0.3200 2.3650 0.5800 ;
        RECT 3.0250 0.3200 3.1150 0.5800 ;
        RECT 4.3500 0.3200 4.4400 0.6050 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 1.2100 1.5500 ;
        RECT 0.0750 1.5500 0.1750 1.8200 ;
        RECT 0.5950 1.5500 0.6950 1.8800 ;
        RECT 1.1100 1.5500 1.2100 1.8800 ;
        RECT 0.0750 0.9500 0.1750 1.4500 ;
        RECT 0.0750 0.8500 1.0100 0.9500 ;
        RECT 0.3900 0.4900 0.4900 0.8500 ;
        RECT 0.9100 0.4900 1.0100 0.8500 ;
    END
    ANTENNADIFFAREA 0.7406 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0450 2.5500 1.1900 ;
        RECT 2.3950 0.8550 2.5500 1.0450 ;
    END
    ANTENNAGATEAREA 0.0576 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1700 1.0500 4.5150 1.1750 ;
    END
    ANTENNAGATEAREA 0.0516 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.5050 3.3500 1.8300 ;
        RECT 3.2500 1.8300 4.2700 1.9200 ;
        RECT 3.0150 1.4250 3.3500 1.5050 ;
        RECT 4.1700 1.5900 4.2700 1.8300 ;
        RECT 3.8100 1.1450 3.9000 1.8300 ;
        RECT 1.7350 1.4150 3.3500 1.4250 ;
        RECT 4.1700 1.4900 4.5400 1.5900 ;
        RECT 3.4250 1.0550 3.9000 1.1450 ;
        RECT 1.7350 1.3250 3.1050 1.4150 ;
        RECT 4.4500 1.3500 4.5400 1.4900 ;
        RECT 3.4250 0.6900 3.5150 1.0550 ;
    END
    ANTENNAGATEAREA 0.1953 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 1.9750 1.8800 2.1450 2.0800 ;
        RECT 0.3400 1.7700 0.4300 2.0800 ;
        RECT 0.8600 1.7700 0.9500 2.0800 ;
        RECT 4.3700 1.7550 4.4600 2.0800 ;
        RECT 2.5250 1.7450 2.6150 2.0800 ;
        RECT 3.0550 1.7450 3.1450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.3000 1.6950 2.4100 1.7850 ;
      RECT 1.3000 0.8100 1.9050 0.9000 ;
      RECT 1.8150 0.4100 1.9050 0.8100 ;
      RECT 1.3000 1.1800 1.3900 1.6950 ;
      RECT 0.5950 1.0900 1.3900 1.1800 ;
      RECT 1.3000 0.9000 1.3900 1.0900 ;
      RECT 2.1600 0.6700 3.1350 0.7600 ;
      RECT 3.0450 0.7600 3.1350 0.8850 ;
      RECT 1.5350 1.2400 1.6250 1.5150 ;
      RECT 1.4800 1.1200 1.6250 1.2400 ;
      RECT 1.4800 1.0300 2.2600 1.1200 ;
      RECT 2.1700 1.1200 2.2600 1.2050 ;
      RECT 2.1600 0.7600 2.2600 1.0300 ;
      RECT 2.7850 1.6050 2.8750 1.9050 ;
      RECT 1.5350 1.5150 2.8750 1.6050 ;
      RECT 2.7650 0.4800 2.8550 0.6700 ;
      RECT 3.6100 1.3250 3.7000 1.7400 ;
      RECT 3.2250 1.2350 3.7000 1.3250 ;
      RECT 3.2250 0.5100 3.6200 0.6000 ;
      RECT 3.5300 0.4100 3.6200 0.5100 ;
      RECT 3.2250 1.1600 3.3150 1.2350 ;
      RECT 2.7850 1.0700 3.3150 1.1600 ;
      RECT 3.2250 0.6000 3.3150 1.0700 ;
      RECT 3.9900 0.7700 4.0800 1.6600 ;
      RECT 3.9100 0.6800 4.0800 0.7700 ;
      RECT 4.6300 1.7450 4.7300 1.9550 ;
      RECT 4.6400 0.9000 4.7300 1.7450 ;
      RECT 4.1700 0.8100 4.7300 0.9000 ;
      RECT 4.6300 0.4100 4.7300 0.8100 ;
      RECT 3.7300 0.5700 3.8200 0.8750 ;
      RECT 3.6300 0.8750 3.8200 0.9650 ;
      RECT 4.1700 0.5700 4.2600 0.8100 ;
      RECT 3.7300 0.4800 4.2600 0.5700 ;
  END
END POSTICG_X5B_A12TH

MACRO POSTICG_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.2500 0.3200 0.3400 0.6000 ;
        RECT 0.7900 0.3200 0.8800 0.6000 ;
        RECT 1.3900 0.3200 1.4800 0.6600 ;
        RECT 2.5500 0.3200 2.7200 0.3400 ;
        RECT 3.7050 0.3200 3.9150 0.5050 ;
        RECT 5.1100 0.3200 5.2000 0.7450 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3350 1.4500 1.4750 1.5500 ;
        RECT 0.3350 1.5500 0.4350 1.8800 ;
        RECT 0.8550 1.5500 0.9550 1.8800 ;
        RECT 1.3750 1.5500 1.4750 1.8800 ;
        RECT 0.4500 0.9500 0.5500 1.4500 ;
        RECT 0.4500 0.8600 1.1800 0.9500 ;
        RECT 0.5050 0.8500 1.1800 0.8600 ;
        RECT 0.5050 0.4550 0.6050 0.8500 ;
        RECT 1.0800 0.4550 1.1800 0.8500 ;
    END
    ANTENNADIFFAREA 0.788 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6400 0.8500 3.7650 1.1900 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.0550 4.9500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0576 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1650 1.2150 2.9850 1.3150 ;
        RECT 2.8950 1.3150 2.9850 1.8300 ;
        RECT 2.1650 1.3150 2.3900 1.3500 ;
        RECT 2.8950 1.8300 3.6150 1.9200 ;
        RECT 3.5250 1.7200 3.6150 1.8300 ;
        RECT 3.5250 1.6300 4.1500 1.7200 ;
        RECT 4.0500 1.7200 4.1500 1.8300 ;
        RECT 4.0500 1.8300 4.9500 1.9200 ;
        RECT 4.8500 1.8000 4.9500 1.8300 ;
        RECT 4.4900 1.2750 4.5800 1.8300 ;
        RECT 4.8500 1.7000 5.3400 1.8000 ;
        RECT 4.2000 1.1850 4.5800 1.2750 ;
        RECT 5.2500 1.2850 5.3400 1.7000 ;
        RECT 4.2000 0.8800 4.2900 1.1850 ;
    END
    ANTENNAGATEAREA 0.2484 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 3.0450 2.0100 3.1350 2.0800 ;
        RECT 5.0500 1.9250 5.1400 2.0800 ;
        RECT 3.7050 1.8400 3.8950 2.0800 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
        RECT 1.1200 1.7700 1.2100 2.0800 ;
        RECT 2.3950 1.7700 2.4850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.5850 0.7200 3.1400 0.8100 ;
      RECT 3.0500 0.5200 3.1400 0.7200 ;
      RECT 2.1350 1.5000 2.7450 1.5900 ;
      RECT 2.6550 1.5900 2.7450 1.9300 ;
      RECT 1.5850 1.1800 1.6750 1.8300 ;
      RECT 0.7550 1.0900 1.6750 1.1800 ;
      RECT 1.5850 0.8100 1.6750 1.0900 ;
      RECT 1.5850 1.8300 2.2250 1.9200 ;
      RECT 2.1350 1.5900 2.2250 1.8300 ;
      RECT 2.0600 0.4300 2.2300 0.7200 ;
      RECT 3.2300 1.3000 3.7700 1.3900 ;
      RECT 3.6800 1.3900 3.7700 1.4250 ;
      RECT 3.6800 1.4250 3.8900 1.5150 ;
      RECT 1.8600 1.0100 1.9500 1.6350 ;
      RECT 3.2300 1.6300 3.4350 1.7200 ;
      RECT 3.2300 1.3900 3.3200 1.6300 ;
      RECT 3.2300 1.0100 3.3200 1.3000 ;
      RECT 1.8600 0.9200 3.3200 1.0100 ;
      RECT 3.2300 0.5000 3.3200 0.9200 ;
      RECT 3.2300 0.4100 3.4350 0.5000 ;
      RECT 4.3100 1.4550 4.4000 1.7200 ;
      RECT 4.0000 1.3650 4.4000 1.4550 ;
      RECT 3.4100 0.6100 4.4000 0.7000 ;
      RECT 4.2300 0.4300 4.4000 0.6100 ;
      RECT 4.0000 0.7000 4.0900 1.3650 ;
      RECT 3.4100 0.7000 3.5000 1.1500 ;
      RECT 4.6700 0.7700 4.7600 1.7200 ;
      RECT 4.6700 0.6800 4.8400 0.7700 ;
      RECT 5.4300 0.9450 5.5200 1.7550 ;
      RECT 4.9300 0.8550 5.5200 0.9450 ;
      RECT 5.4300 0.6050 5.5200 0.8550 ;
      RECT 4.4900 0.5700 4.5800 1.0750 ;
      RECT 4.9300 0.5700 5.0200 0.8550 ;
      RECT 4.4900 0.4800 5.0200 0.5700 ;
  END
END POSTICG_X6B_A12TH

MACRO POSTICG_X7P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 1.0700 0.3200 1.1600 0.6500 ;
        RECT 1.6250 0.3200 1.7150 0.6500 ;
        RECT 2.2400 0.3200 2.3300 0.6000 ;
        RECT 3.2350 0.3200 3.3250 0.6000 ;
        RECT 4.4400 0.3200 4.5300 0.4100 ;
        RECT 5.9050 0.3200 5.9950 0.5000 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3300 1.2450 2.0000 1.3550 ;
        RECT 0.3300 1.3550 0.4400 1.7600 ;
        RECT 0.8500 1.3550 0.9600 1.7600 ;
        RECT 1.3700 1.3550 1.4800 1.7600 ;
        RECT 1.8900 1.3550 2.0000 1.7600 ;
        RECT 0.4450 0.9550 0.5550 1.2450 ;
        RECT 0.4450 0.8450 2.0000 0.9550 ;
        RECT 0.7800 0.4700 0.8900 0.8450 ;
        RECT 1.3400 0.4700 1.4500 0.8450 ;
        RECT 1.8900 0.4700 2.0000 0.8450 ;
    END
    ANTENNADIFFAREA 1.0472 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.8100 4.5500 1.0100 ;
        RECT 4.3550 1.0100 4.5500 1.1250 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7350 0.9800 5.9500 1.1900 ;
        RECT 5.8450 0.8950 5.9500 0.9800 ;
    END
    ANTENNAGATEAREA 0.0669 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5800 1.2950 2.9500 1.3500 ;
        RECT 2.5800 1.1950 3.7500 1.2950 ;
        RECT 3.6500 1.2950 3.7500 1.7900 ;
        RECT 2.5800 1.1850 2.9500 1.1950 ;
        RECT 3.6500 1.7900 4.4850 1.8800 ;
        RECT 4.3950 1.5500 4.4850 1.7900 ;
        RECT 4.3950 1.4600 4.9650 1.5500 ;
        RECT 4.8750 1.5500 4.9650 1.8300 ;
        RECT 4.8750 1.8300 5.8450 1.9200 ;
        RECT 5.7550 1.5900 5.8450 1.8300 ;
        RECT 5.3450 1.3300 5.4350 1.8300 ;
        RECT 5.7550 1.5000 6.1400 1.5900 ;
        RECT 5.3450 1.1900 5.4550 1.3300 ;
        RECT 6.0500 1.1550 6.1400 1.5000 ;
        RECT 5.0850 1.1000 5.4550 1.1900 ;
        RECT 5.0850 1.0800 5.1750 1.1000 ;
        RECT 4.9550 0.9900 5.1750 1.0800 ;
        RECT 4.9550 0.8700 5.0450 0.9900 ;
    END
    ANTENNAGATEAREA 0.3033 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 3.5400 2.0250 3.9500 2.0800 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 0.6000 1.7500 0.6900 2.0800 ;
        RECT 1.1200 1.7500 1.2100 2.0800 ;
        RECT 1.6400 1.7500 1.7300 2.0800 ;
        RECT 2.1600 1.7500 2.2500 2.0800 ;
        RECT 2.9100 1.7500 3.0000 2.0800 ;
        RECT 5.9350 1.7100 6.0250 2.0800 ;
        RECT 4.5750 1.6800 4.7450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1600 0.6900 3.7850 0.7800 ;
      RECT 3.6950 0.4100 3.7850 0.6900 ;
      RECT 2.1600 1.4550 3.2900 1.5450 ;
      RECT 3.2000 1.5450 3.2900 1.9500 ;
      RECT 2.1600 1.1400 2.2500 1.4550 ;
      RECT 0.7000 1.0500 2.2500 1.1400 ;
      RECT 2.1600 0.7800 2.2500 1.0500 ;
      RECT 2.6200 1.5450 2.7100 1.9400 ;
      RECT 2.7250 0.4100 2.8150 0.6900 ;
      RECT 2.3400 0.9600 2.4300 1.1900 ;
      RECT 2.3400 0.8700 3.9750 0.9600 ;
      RECT 3.8850 0.7600 4.0700 0.8500 ;
      RECT 3.8850 0.8500 3.9750 0.8700 ;
      RECT 3.8850 1.2600 4.6850 1.3500 ;
      RECT 3.8850 0.9600 3.9750 1.2600 ;
      RECT 3.9800 0.4300 4.0700 0.7600 ;
      RECT 4.1300 1.5900 4.3050 1.6800 ;
      RECT 4.2150 1.3500 4.3050 1.5900 ;
      RECT 3.1000 0.8700 3.4700 1.1050 ;
      RECT 5.1350 1.3700 5.2250 1.7400 ;
      RECT 4.7750 1.2800 5.2250 1.3700 ;
      RECT 4.1700 0.6100 5.1750 0.7000 ;
      RECT 5.0850 0.7000 5.1750 0.7800 ;
      RECT 5.0850 0.4100 5.1750 0.6100 ;
      RECT 4.7750 0.7000 4.8650 1.2800 ;
      RECT 4.1700 0.7000 4.2600 0.9800 ;
      RECT 4.0650 0.9800 4.2600 1.0700 ;
      RECT 5.5450 0.7700 5.6350 1.7400 ;
      RECT 5.4650 0.6800 5.6350 0.7700 ;
      RECT 6.2300 0.7000 6.3200 1.9000 ;
      RECT 5.7250 0.6100 6.3200 0.7000 ;
      RECT 5.2850 0.5700 5.3750 1.0100 ;
      RECT 5.7250 0.5700 5.8150 0.6100 ;
      RECT 5.2850 0.4800 5.8150 0.5700 ;
  END
END POSTICG_X7P5B_A12TH

MACRO POSTICG_X9B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6000 ;
        RECT 0.6000 0.3200 0.6900 0.6000 ;
        RECT 1.1200 0.3200 1.2100 0.6000 ;
        RECT 1.6400 0.3200 1.7300 0.6000 ;
        RECT 2.6850 0.3200 2.8550 0.3650 ;
        RECT 3.7800 0.3200 3.8700 0.5800 ;
        RECT 4.6450 0.3200 4.7350 0.5800 ;
        RECT 5.8950 0.3200 6.0650 0.3600 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4350 2.0350 1.5650 ;
        RECT 1.9050 1.5650 2.0350 1.6600 ;
        RECT 0.0800 1.5650 0.1700 1.8300 ;
        RECT 0.6000 1.5650 0.6900 1.8300 ;
        RECT 1.1200 1.5650 1.2100 1.8300 ;
        RECT 1.6400 1.5650 1.7300 1.8300 ;
        RECT 0.2500 0.9500 0.3650 1.4350 ;
        RECT 1.9050 1.6600 2.2500 1.7900 ;
        RECT 0.2500 0.8200 1.4700 0.9500 ;
        RECT 2.1600 1.7900 2.2500 1.9200 ;
        RECT 0.3400 0.4750 0.4300 0.8200 ;
        RECT 0.8600 0.4750 0.9500 0.8200 ;
        RECT 1.3800 0.4600 1.4700 0.8200 ;
    END
    ANTENNADIFFAREA 1.2012 ;
  END ECK

  PIN SEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7800 1.0500 4.2000 1.1500 ;
    END
    ANTENNAGATEAREA 0.0888 ;
  END SEN

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.9500 5.9500 1.1900 ;
        RECT 5.8500 0.8500 6.1550 0.9500 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3450 1.2800 3.7500 1.3750 ;
        RECT 3.6500 1.3750 3.7500 1.6400 ;
        RECT 2.3450 1.2750 3.4600 1.2800 ;
        RECT 3.6500 1.6400 5.1450 1.7300 ;
        RECT 3.2100 1.2000 3.4600 1.2750 ;
        RECT 2.3450 0.9900 2.4350 1.2750 ;
        RECT 5.0550 1.7300 5.1450 1.8300 ;
        RECT 2.2500 0.9000 2.4350 0.9900 ;
        RECT 5.0550 1.8300 6.0900 1.9200 ;
        RECT 6.0000 1.3900 6.0900 1.8300 ;
        RECT 5.4500 1.2100 5.5400 1.8300 ;
        RECT 6.0000 1.2800 6.1750 1.3900 ;
        RECT 5.0450 1.1200 5.5400 1.2100 ;
        RECT 5.0450 0.7150 5.1350 1.1200 ;
    END
    ANTENNAGATEAREA 0.3576 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 5.9100 2.0100 6.0000 2.0800 ;
        RECT 3.8400 1.9300 3.9300 2.0800 ;
        RECT 1.8600 1.8800 2.0300 2.0800 ;
        RECT 4.4950 1.8700 4.8650 2.0800 ;
        RECT 3.1600 1.8400 3.2500 2.0800 ;
        RECT 0.3400 1.7700 0.4300 2.0800 ;
        RECT 0.8600 1.7700 0.9500 2.0800 ;
        RECT 1.3800 1.7700 1.4700 2.0800 ;
        RECT 2.4200 1.7700 2.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1450 1.4800 3.5100 1.5700 ;
      RECT 3.4200 1.5700 3.5100 1.9100 ;
      RECT 3.0300 0.8650 3.2900 0.9550 ;
      RECT 3.2000 0.6600 3.2900 0.8650 ;
      RECT 2.1450 1.2200 2.2350 1.4800 ;
      RECT 0.9000 1.1300 2.2350 1.2200 ;
      RECT 2.0500 0.8100 2.1400 1.1300 ;
      RECT 2.1900 0.6600 2.4000 0.7200 ;
      RECT 2.9000 1.5700 2.9900 1.9100 ;
      RECT 2.0500 0.7200 2.6150 0.8100 ;
      RECT 2.5250 0.8100 2.6150 1.0900 ;
      RECT 2.5250 1.0900 3.1200 1.1800 ;
      RECT 3.0300 0.9550 3.1200 1.0900 ;
      RECT 4.3000 0.7600 4.7550 0.7800 ;
      RECT 4.6650 0.7800 4.7550 0.8800 ;
      RECT 3.5200 0.6700 4.7550 0.7600 ;
      RECT 3.5900 0.7600 3.6800 1.1000 ;
      RECT 1.8500 0.5700 1.9400 1.0400 ;
      RECT 2.8500 0.5700 2.9400 0.9100 ;
      RECT 2.7250 0.9100 2.9400 1.0000 ;
      RECT 3.5200 0.5700 3.6100 0.6700 ;
      RECT 1.8500 0.4800 3.6100 0.5700 ;
      RECT 4.1000 1.4400 4.3900 1.5300 ;
      RECT 4.3000 0.7800 4.3900 1.4400 ;
      RECT 4.4150 0.4100 4.5050 0.6700 ;
      RECT 5.2700 1.4400 5.3600 1.6800 ;
      RECT 4.8450 1.3500 5.3600 1.4400 ;
      RECT 4.8450 0.4800 5.3200 0.5700 ;
      RECT 5.2300 0.5700 5.3200 0.6950 ;
      RECT 4.8450 1.2500 4.9350 1.3500 ;
      RECT 4.4950 1.1600 4.9350 1.2500 ;
      RECT 4.8450 0.5700 4.9350 1.1600 ;
      RECT 4.4950 1.0400 4.5850 1.1600 ;
      RECT 5.6300 0.7500 5.7200 1.6700 ;
      RECT 5.6300 0.6600 5.8250 0.7500 ;
      RECT 6.2300 1.5500 6.3200 1.6700 ;
      RECT 6.2300 1.4650 6.3550 1.5500 ;
      RECT 6.2650 0.7450 6.3550 1.4650 ;
      RECT 6.2300 0.6550 6.3550 0.7450 ;
      RECT 5.9350 0.5700 6.3550 0.6550 ;
      RECT 5.4300 0.5650 6.3550 0.5700 ;
      RECT 5.4300 0.4800 6.0250 0.5650 ;
      RECT 5.4300 0.5700 5.5200 0.8950 ;
      RECT 5.3150 0.8950 5.5200 0.9850 ;
  END
END POSTICG_X9B_A12TH

MACRO PREICG_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5450 ;
        RECT 0.5950 0.3200 0.6950 0.5700 ;
        RECT 2.0100 0.3200 2.1000 0.8050 ;
        RECT 2.9450 0.3200 3.0450 0.5100 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.1000 0.7500 1.5000 ;
        RECT 0.6500 1.5000 0.8900 1.6000 ;
        RECT 0.6500 1.0000 0.9050 1.1000 ;
        RECT 0.7900 1.6000 0.8900 1.8200 ;
        RECT 0.7900 1.8200 2.1250 1.9200 ;
        RECT 2.0250 1.4150 2.1250 1.8200 ;
        RECT 2.0250 1.3150 2.7200 1.4150 ;
        RECT 2.6200 1.1950 2.7200 1.3150 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7000 0.1650 1.1550 ;
    END
    ANTENNAGATEAREA 0.0282 ;
  END E

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.5200 3.3500 1.6200 ;
        RECT 3.2300 1.6200 3.3500 1.9900 ;
        RECT 3.1600 0.4200 3.3500 0.5200 ;
    END
    ANTENNADIFFAREA 0.11105 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 2.9300 1.9600 3.0300 2.0800 ;
        RECT 2.4200 1.8700 2.5150 2.0800 ;
        RECT 0.5950 1.7800 0.6950 2.0800 ;
        RECT 2.2350 1.5050 2.3300 2.0800 ;
        RECT 2.9300 1.8650 3.1200 1.9600 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.2450 0.5500 1.6850 ;
    END
    ANTENNAGATEAREA 0.0363 ;
  END SE
  OBS
    LAYER M1 ;
      RECT 1.2050 1.4450 1.3750 1.5500 ;
      RECT 0.9950 1.3550 1.3750 1.4450 ;
      RECT 0.9950 0.8350 1.0850 1.3550 ;
      RECT 0.2600 0.7600 1.0850 0.8350 ;
      RECT 0.2600 0.7450 1.2000 0.7600 ;
      RECT 0.9950 0.6700 1.2000 0.7450 ;
      RECT 0.2600 0.4400 0.4800 0.5300 ;
      RECT 0.2600 0.8350 0.3500 1.3000 ;
      RECT 0.0500 1.3000 0.3500 1.3900 ;
      RECT 0.2600 0.5300 0.3500 0.7450 ;
      RECT 0.0500 1.3900 0.1700 1.8900 ;
      RECT 0.9800 1.6400 1.5550 1.7300 ;
      RECT 0.9800 1.5550 1.0700 1.6400 ;
      RECT 1.4650 1.2650 1.5550 1.6400 ;
      RECT 1.3100 1.1750 1.7450 1.2650 ;
      RECT 1.3100 1.0600 1.4000 1.1750 ;
      RECT 1.1750 0.8900 1.4000 1.0600 ;
      RECT 1.3100 0.5700 1.4000 0.8900 ;
      RECT 0.8450 0.4800 1.4000 0.5700 ;
      RECT 0.8450 0.4200 1.0150 0.4800 ;
      RECT 1.4900 0.9450 2.3000 1.0350 ;
      RECT 2.2100 0.8350 2.3000 0.9450 ;
      RECT 1.6650 1.5250 1.7550 1.6350 ;
      RECT 1.6650 1.4350 1.9350 1.5250 ;
      RECT 1.8450 1.0350 1.9350 1.4350 ;
      RECT 1.4900 0.6250 1.5800 0.9450 ;
      RECT 2.4400 1.5050 2.9200 1.5950 ;
      RECT 2.8200 0.9950 2.9200 1.5050 ;
      RECT 2.4100 0.9050 2.9200 0.9950 ;
      RECT 2.4100 0.9950 2.5000 1.1350 ;
      RECT 2.4100 0.7450 2.5000 0.9050 ;
      RECT 2.0700 1.1350 2.5000 1.2250 ;
      RECT 2.2250 0.6550 2.5000 0.7450 ;
      RECT 2.7400 1.6850 3.1400 1.7750 ;
      RECT 3.0500 1.3950 3.1400 1.6850 ;
      RECT 3.0500 1.0050 3.1600 1.3950 ;
      RECT 3.0500 0.7300 3.1400 1.0050 ;
      RECT 2.5900 0.6400 3.1400 0.7300 ;
      RECT 2.6200 1.8700 2.8300 1.9600 ;
      RECT 2.7400 1.7750 2.8300 1.8700 ;
      RECT 2.5900 0.5150 2.6800 0.6400 ;
      RECT 2.3600 0.4250 2.6800 0.5150 ;
  END
END PREICG_X0P5B_A12TH

MACRO OR2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.5150 0.3200 0.6050 0.8600 ;
        RECT 1.1100 0.3200 1.2000 0.6350 ;
        RECT 1.6300 0.3200 1.7200 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.0500 0.8200 1.1500 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1300 1.2500 1.0300 1.3500 ;
        RECT 0.9300 1.0200 1.0300 1.2500 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3650 1.2500 1.7500 1.3500 ;
        RECT 1.3650 1.3500 1.4650 1.7200 ;
        RECT 1.6500 0.9500 1.7500 1.2500 ;
        RECT 1.3650 0.8500 1.7500 0.9500 ;
        RECT 1.3650 0.4900 1.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.6300 1.8400 1.7200 2.0800 ;
        RECT 1.0950 1.7700 1.1850 2.0800 ;
        RECT 0.1350 1.7000 0.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1400 1.0550 1.5300 1.1450 ;
      RECT 0.5850 1.5000 1.2300 1.5900 ;
      RECT 1.1400 1.1450 1.2300 1.5000 ;
      RECT 1.1400 0.9000 1.2300 1.0550 ;
      RECT 0.7750 0.8100 1.2300 0.9000 ;
      RECT 0.5850 1.5900 0.6750 1.9300 ;
      RECT 0.7750 0.4900 0.8650 0.8100 ;
  END
END OR2_X2M_A12TH

MACRO OR2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.5150 0.3200 0.6050 0.6500 ;
        RECT 1.0500 0.3200 1.1400 0.6500 ;
        RECT 1.5700 0.3200 1.6600 0.6500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1850 1.2500 1.0250 1.3500 ;
        RECT 0.1850 1.1550 0.2750 1.2500 ;
        RECT 0.9250 1.0000 1.0250 1.2500 ;
        RECT 0.0750 1.0500 0.2750 1.1550 ;
    END
    ANTENNAGATEAREA 0.1476 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3850 1.0500 0.8050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1476 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3050 1.2500 1.9500 1.3500 ;
        RECT 1.3050 1.3500 1.4050 1.7200 ;
        RECT 1.8300 1.3500 1.9500 1.7200 ;
        RECT 1.8500 0.9500 1.9500 1.2500 ;
        RECT 1.3050 0.8500 1.9500 0.9500 ;
        RECT 1.3050 0.5050 1.4050 0.8500 ;
        RECT 1.8300 0.5050 1.9500 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.5700 1.8400 1.6600 2.0800 ;
        RECT 1.0500 1.7400 1.1400 2.0800 ;
        RECT 0.0800 1.7300 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1200 1.0550 1.6250 1.1450 ;
      RECT 0.5300 1.5900 0.6200 1.9300 ;
      RECT 0.7750 0.4600 0.8650 0.8000 ;
      RECT 0.5300 1.5000 1.2100 1.5900 ;
      RECT 1.1200 1.1450 1.2100 1.5000 ;
      RECT 1.1200 0.8900 1.2100 1.0550 ;
      RECT 0.7750 0.8000 1.2100 0.8900 ;
  END
END OR2_X3M_A12TH

MACRO OR2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.4600 0.3200 0.5500 0.7200 ;
        RECT 0.9800 0.3200 1.0700 0.6950 ;
        RECT 1.5750 0.3200 1.6650 0.6250 ;
        RECT 2.0950 0.3200 2.1850 0.6250 ;
        RECT 2.6150 0.3200 2.7050 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.2500 1.4200 1.3500 ;
        RECT 0.4100 1.1600 0.7350 1.2500 ;
        RECT 1.3200 1.0000 1.4200 1.2500 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.0700 1.2100 1.1500 ;
        RECT 0.2400 0.9700 1.2100 1.0700 ;
        RECT 0.2400 0.8550 0.3500 0.9700 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8300 1.2500 2.5500 1.3500 ;
        RECT 1.8300 1.3500 1.9300 1.7200 ;
        RECT 2.3500 1.3500 2.4500 1.7200 ;
        RECT 2.4500 0.9500 2.5500 1.2500 ;
        RECT 1.8300 0.8500 2.5500 0.9500 ;
        RECT 1.8300 0.4850 1.9300 0.8500 ;
        RECT 2.3500 0.4850 2.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.0950 1.8400 2.1850 2.0800 ;
        RECT 2.6150 1.8400 2.7050 2.0800 ;
        RECT 0.5300 1.7300 0.6200 2.0800 ;
        RECT 1.5000 1.7300 1.5900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.5300 1.0550 2.2200 1.1450 ;
      RECT 0.0800 1.5900 0.1700 1.9300 ;
      RECT 0.7150 0.4400 0.8150 0.7900 ;
      RECT 1.2350 0.4400 1.3350 0.7900 ;
      RECT 0.9800 1.5900 1.0700 1.8700 ;
      RECT 0.0800 1.5000 1.6200 1.5900 ;
      RECT 1.5300 1.1450 1.6200 1.5000 ;
      RECT 1.5300 0.8800 1.6200 1.0550 ;
      RECT 0.7150 0.7900 1.6200 0.8800 ;
  END
END OR2_X4M_A12TH

MACRO OR2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.5900 ;
        RECT 2.7050 0.3200 2.8050 0.6350 ;
        RECT 3.2250 0.3200 3.3250 0.6350 ;
        RECT 3.7500 0.3200 3.8500 0.6350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.9500 3.3500 1.2500 ;
        RECT 2.4450 1.2500 3.5850 1.3500 ;
        RECT 2.4450 0.8500 3.5850 0.9500 ;
        RECT 2.4450 1.3500 2.5450 1.7350 ;
        RECT 2.9650 1.3500 3.0650 1.7350 ;
        RECT 3.4850 1.3500 3.5850 1.7350 ;
        RECT 2.4450 0.4900 2.5450 0.8500 ;
        RECT 2.9650 0.4900 3.0650 0.8500 ;
        RECT 3.4850 0.4900 3.5850 0.8500 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0500 2.1150 1.1500 ;
        RECT 2.0150 0.7250 2.1150 1.0500 ;
        RECT 0.2450 0.7200 0.3450 1.0500 ;
    END
    ANTENNAGATEAREA 0.2988 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 0.8500 1.8900 0.9500 ;
    END
    ANTENNAGATEAREA 0.2988 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 2.1800 1.7700 2.2800 2.0800 ;
        RECT 2.7050 1.7700 2.8050 2.0800 ;
        RECT 3.2250 1.7700 3.3250 2.0800 ;
        RECT 3.7500 1.7700 3.8500 2.0800 ;
        RECT 0.0900 1.7250 0.1900 2.0800 ;
        RECT 1.1300 1.7250 1.2300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2350 1.0600 3.0750 1.1500 ;
      RECT 0.6100 1.5650 0.7100 1.9050 ;
      RECT 0.3150 0.4350 0.4850 0.5200 ;
      RECT 0.8350 0.4350 1.0050 0.5200 ;
      RECT 1.8750 0.4350 2.0450 0.5200 ;
      RECT 1.6500 1.5650 1.7500 1.9050 ;
      RECT 1.3550 0.4350 1.5250 0.5200 ;
      RECT 0.6100 1.4750 2.3250 1.5650 ;
      RECT 2.2350 1.1500 2.3250 1.4750 ;
      RECT 2.2350 0.6950 2.3250 1.0600 ;
      RECT 2.2350 0.6100 2.3400 0.6950 ;
      RECT 0.3150 0.5200 2.3400 0.6100 ;
  END
END OR2_X6M_A12TH

MACRO OR2_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 1.3150 0.3200 1.4050 0.6500 ;
        RECT 1.7950 0.3200 1.9650 0.5500 ;
        RECT 2.3150 0.3200 2.4850 0.5500 ;
        RECT 2.9100 0.3200 3.0800 0.5500 ;
        RECT 3.4700 0.3200 3.5600 0.6500 ;
        RECT 3.9900 0.3200 4.0800 0.6500 ;
        RECT 4.5100 0.3200 4.6000 0.6500 ;
        RECT 5.0300 0.3200 5.1200 0.6500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9100 0.8500 2.8750 0.9300 ;
        RECT 0.4750 0.9300 2.8750 0.9500 ;
        RECT 0.4750 0.9500 1.0100 1.0400 ;
        RECT 1.7400 0.9500 2.1100 1.0600 ;
        RECT 2.7650 0.9500 2.8750 1.1700 ;
    END
    ANTENNAGATEAREA 0.4032 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.2900 2.3400 1.3500 ;
        RECT 0.6950 1.2600 2.6300 1.2900 ;
        RECT 0.3850 1.2500 2.6300 1.2600 ;
        RECT 1.4000 1.1800 1.6100 1.2500 ;
        RECT 2.2200 1.1750 2.6300 1.2500 ;
        RECT 0.3850 1.1600 0.7950 1.2500 ;
    END
    ANTENNAGATEAREA 0.4032 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2050 1.4350 4.9650 1.5650 ;
        RECT 3.2050 1.5650 3.3050 1.9200 ;
        RECT 3.7250 1.5650 3.8250 1.9200 ;
        RECT 4.2450 1.5650 4.3450 1.9200 ;
        RECT 4.7650 1.5650 4.8650 1.9200 ;
        RECT 4.8350 0.9650 4.9650 1.4350 ;
        RECT 3.2050 0.8350 4.9650 0.9650 ;
        RECT 3.2050 0.5050 3.3050 0.8350 ;
        RECT 3.7250 0.5050 3.8250 0.8350 ;
        RECT 4.2450 0.5050 4.3450 0.8350 ;
        RECT 4.7650 0.5050 4.8650 0.8350 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 3.4700 1.7700 3.5600 2.0800 ;
        RECT 3.9900 1.7700 4.0800 2.0800 ;
        RECT 4.5100 1.7700 4.6000 2.0800 ;
        RECT 5.0300 1.7700 5.1200 2.0800 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 1.0100 1.7500 1.1000 2.0800 ;
        RECT 1.9100 1.7500 2.0000 2.0800 ;
        RECT 2.9500 1.7500 3.0400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.9950 1.0700 4.7000 1.1600 ;
      RECT 0.5600 1.5900 0.6500 1.9300 ;
      RECT 1.4600 1.5900 1.5500 1.9400 ;
      RECT 1.5350 0.4100 1.7050 0.6700 ;
      RECT 2.0950 0.4100 2.1850 0.6700 ;
      RECT 2.4150 1.5900 2.5050 1.9300 ;
      RECT 2.6150 0.4100 2.7050 0.6700 ;
      RECT 0.5600 1.5000 3.0850 1.5900 ;
      RECT 2.9950 1.1600 3.0850 1.5000 ;
      RECT 2.9950 0.7600 3.0850 1.0700 ;
      RECT 1.5350 0.6700 3.0850 0.7600 ;
  END
END OR2_X8M_A12TH

MACRO OR3_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.5200 ;
        RECT 0.8650 0.3200 1.0350 0.5200 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 0.8100 0.3500 1.1600 ;
    END
    ANTENNAGATEAREA 0.0531 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.8050 0.5600 1.3000 ;
    END
    ANTENNAGATEAREA 0.0531 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.5650 1.3500 1.3150 ;
        RECT 1.1750 1.3150 1.3500 1.4150 ;
        RECT 1.1400 0.4650 1.3500 0.5650 ;
        RECT 1.1750 1.4150 1.2750 1.7600 ;
    END
    ANTENNADIFFAREA 0.167075 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9150 1.3800 1.0150 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.8400 1.1000 ;
    END
    ANTENNAGATEAREA 0.0531 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.0500 0.6100 1.0500 0.7000 ;
      RECT 0.9600 0.7000 1.0500 0.7100 ;
      RECT 0.9600 0.7100 1.1000 0.9000 ;
      RECT 0.0850 1.7900 0.2550 1.9900 ;
      RECT 0.0500 1.7000 0.2550 1.7900 ;
      RECT 0.0500 0.7000 0.1400 1.7000 ;
      RECT 0.1250 0.4200 0.2150 0.6100 ;
      RECT 0.6450 0.4150 0.7350 0.6100 ;
  END
END OR3_X0P5M_A12TH

MACRO OR3_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.7200 ;
        RECT 0.8650 0.3200 1.0350 0.7200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.8800 1.6400 1.0500 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0100 0.8400 1.3900 ;
    END
    ANTENNAGATEAREA 0.0669 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0100 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0669 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0100 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0669 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8000 1.3500 1.3150 ;
        RECT 1.1750 1.3150 1.3500 1.4150 ;
        RECT 1.1750 0.7000 1.3500 0.8000 ;
        RECT 1.1750 1.4150 1.2750 1.7600 ;
        RECT 1.1750 0.4150 1.2750 0.7000 ;
    END
    ANTENNADIFFAREA 0.236775 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0500 0.8100 1.0500 0.9000 ;
      RECT 0.9600 0.9000 1.0500 0.9300 ;
      RECT 0.9600 0.9300 1.1000 1.1000 ;
      RECT 0.0850 1.7900 0.2550 1.9900 ;
      RECT 0.0500 1.7000 0.2550 1.7900 ;
      RECT 0.0500 0.9000 0.1400 1.7000 ;
      RECT 0.1250 0.6100 0.2150 0.8100 ;
      RECT 0.6450 0.5900 0.7350 0.8100 ;
  END
END OR3_X0P7M_A12TH

MACRO OR3_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.7850 0.3200 0.8750 0.5700 ;
        RECT 1.3300 0.3200 1.5000 0.5350 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0850 0.8400 1.3050 0.9500 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3650 1.0500 1.1150 1.1600 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8050 1.4500 1.1000 1.5500 ;
        RECT 0.8050 1.4200 0.9650 1.4500 ;
        RECT 0.5550 1.3250 0.9650 1.4200 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9050 1.7500 1.2900 ;
        RECT 1.6300 1.2900 1.7500 1.7200 ;
        RECT 1.6300 0.4950 1.7500 0.9050 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.3300 1.8350 1.5000 2.0800 ;
        RECT 0.0800 1.7300 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6800 1.6500 1.5400 1.7400 ;
      RECT 1.4500 0.7500 1.5400 1.6500 ;
      RECT 0.5250 0.6600 1.5400 0.7500 ;
      RECT 0.5250 0.5200 0.6150 0.6600 ;
      RECT 0.6800 1.7400 0.8500 1.9600 ;
      RECT 1.0450 0.5200 1.1350 0.6600 ;
  END
END OR3_X1M_A12TH

MACRO OR3_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.6350 ;
        RECT 0.6400 0.3200 0.7400 0.5100 ;
        RECT 1.1500 0.3200 1.3200 0.5700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.2500 ;
        RECT 0.0500 1.2500 0.4800 1.3500 ;
        RECT 0.0500 0.8500 0.4800 0.9500 ;
        RECT 0.3800 1.3500 0.4800 1.8100 ;
        RECT 0.3800 0.5050 0.4800 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9800 0.8500 1.8800 0.9500 ;
    END
    ANTENNAGATEAREA 0.1254 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 2.0200 1.3500 ;
        RECT 0.7700 1.1050 0.8700 1.2500 ;
        RECT 1.9200 1.0950 2.0200 1.2500 ;
    END
    ANTENNAGATEAREA 0.1254 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2050 1.0500 1.6950 1.1500 ;
    END
    ANTENNAGATEAREA 0.1254 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 2.0250 1.7700 2.1250 2.0800 ;
        RECT 0.6550 1.6450 0.7550 2.0800 ;
        RECT 0.1200 1.5950 0.2200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.3700 1.5450 1.4600 1.8900 ;
      RECT 0.5800 1.4550 1.4600 1.5450 ;
      RECT 0.5800 0.6600 1.5900 0.7500 ;
      RECT 1.4200 0.4100 1.5900 0.6600 ;
      RECT 0.8900 0.4100 1.0600 0.6600 ;
      RECT 0.5800 1.1500 0.6700 1.4550 ;
      RECT 0.3250 1.0600 0.6700 1.1500 ;
      RECT 0.5800 0.7500 0.6700 1.0600 ;
  END
END OR3_X1P4M_A12TH

MACRO OR3_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6550 ;
        RECT 0.6350 0.3200 0.8050 0.5450 ;
        RECT 1.9450 0.3200 2.1150 0.5450 ;
        RECT 2.6250 0.3200 2.7250 0.6050 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1800 0.8500 1.3800 0.9500 ;
        RECT 1.2800 0.9500 1.3800 1.0300 ;
        RECT 0.1800 0.9500 0.2800 1.3400 ;
        RECT 1.2800 1.0300 1.5900 1.1300 ;
    END
    ANTENNAGATEAREA 0.1719 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0900 1.2500 1.8650 1.3500 ;
        RECT 1.7750 1.1650 1.8650 1.2500 ;
        RECT 1.0900 1.1400 1.1900 1.2500 ;
        RECT 0.7200 1.0400 1.1900 1.1400 ;
    END
    ANTENNAGATEAREA 0.1719 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.2500 0.9700 1.3700 ;
        RECT 0.8700 1.3700 0.9700 1.4500 ;
        RECT 0.8700 1.4500 2.0750 1.5500 ;
        RECT 1.9750 1.0400 2.0750 1.4500 ;
        RECT 1.7950 0.9400 2.0750 1.0400 ;
    END
    ANTENNAGATEAREA 0.1719 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9500 2.7500 1.2500 ;
        RECT 2.3650 1.2500 2.7500 1.3500 ;
        RECT 2.3650 0.8500 2.7500 0.9500 ;
        RECT 2.3650 1.3500 2.4650 1.7250 ;
        RECT 2.3650 0.5050 2.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.7200 1.8750 0.8900 2.0800 ;
        RECT 2.0700 1.8750 2.2400 2.0800 ;
        RECT 2.6250 1.7700 2.7250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1700 1.0450 2.5250 1.1450 ;
      RECT 0.0750 1.6500 2.2700 1.7500 ;
      RECT 2.1700 1.1450 2.2700 1.6500 ;
      RECT 2.1700 0.7500 2.2700 1.0450 ;
      RECT 0.3700 0.6500 2.2700 0.7500 ;
      RECT 0.0750 1.7500 0.1750 1.9100 ;
      RECT 0.0750 1.4950 0.1750 1.6500 ;
      RECT 0.3700 0.5400 0.4700 0.6500 ;
      RECT 1.6050 0.4550 1.7750 0.6500 ;
      RECT 1.3800 1.7500 1.5500 1.9400 ;
  END
END OR3_X2M_A12TH

MACRO OR3_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 1.1300 0.3200 1.3000 0.6250 ;
        RECT 1.7750 0.3200 1.8750 0.4800 ;
        RECT 2.3150 0.3200 2.4150 0.4800 ;
        RECT 2.8400 0.3200 2.9400 0.4800 ;
        RECT 3.3600 0.3200 3.4700 0.6050 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6000 0.8500 2.5650 0.9100 ;
        RECT 1.7750 0.9100 2.5650 0.9500 ;
        RECT 0.6000 0.8100 1.9100 0.8500 ;
        RECT 2.4500 0.9500 2.5650 1.1300 ;
        RECT 0.6000 0.7650 1.0150 0.8100 ;
    END
    ANTENNAGATEAREA 0.252 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6750 1.0500 2.2950 1.1100 ;
        RECT 1.5800 1.1100 2.2950 1.1500 ;
        RECT 0.6750 1.0100 1.6700 1.0500 ;
    END
    ANTENNAGATEAREA 0.252 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1800 1.2500 2.8300 1.3500 ;
        RECT 1.2550 1.2100 1.4750 1.2500 ;
        RECT 0.1800 1.0600 0.2800 1.2500 ;
        RECT 2.7300 0.9850 2.8300 1.2500 ;
    END
    ANTENNAGATEAREA 0.252 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1050 0.8500 3.7450 0.9500 ;
        RECT 3.6450 0.9500 3.7450 1.2700 ;
        RECT 3.6300 0.5500 3.7450 0.8500 ;
        RECT 3.1050 0.5350 3.2050 0.8500 ;
        RECT 3.1050 1.2700 3.7450 1.3700 ;
        RECT 3.1050 1.3700 3.2050 1.7150 ;
        RECT 3.6300 1.3700 3.7450 1.7100 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.0750 1.8050 0.1750 2.0800 ;
        RECT 1.3950 1.8050 1.4950 2.0800 ;
        RECT 3.3650 1.7900 3.4650 2.0800 ;
        RECT 2.8400 1.7600 2.9400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.9250 1.0700 3.4100 1.1600 ;
      RECT 0.7350 1.6000 0.8350 1.9500 ;
      RECT 2.0550 1.6000 2.1550 1.9550 ;
      RECT 0.7350 1.5100 3.0150 1.6000 ;
      RECT 2.9250 1.1600 3.0150 1.5100 ;
      RECT 2.9250 0.6800 3.0150 1.0700 ;
      RECT 1.4350 0.5900 3.0150 0.6800 ;
  END
END OR3_X3M_A12TH

MACRO OR3_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 2.0700 0.3200 2.1700 0.4350 ;
        RECT 2.5900 0.3200 2.6900 0.5800 ;
        RECT 3.1100 0.3200 3.2100 0.5800 ;
        RECT 3.6350 0.3200 3.7350 0.5800 ;
        RECT 4.1550 0.3200 4.2550 0.6400 ;
        RECT 4.6750 0.3200 4.7750 0.6400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9000 1.0500 4.5100 1.1500 ;
        RECT 3.9000 1.1500 3.9900 1.6350 ;
        RECT 4.4200 1.1500 4.5100 1.6350 ;
        RECT 3.9000 0.5500 3.9900 1.0500 ;
        RECT 4.4200 0.5500 4.5100 1.0500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7000 0.8500 3.5650 0.9500 ;
        RECT 1.9950 0.9500 3.5650 0.9600 ;
        RECT 1.7000 0.7600 1.8000 0.8500 ;
        RECT 1.9950 0.9600 2.2000 1.0100 ;
        RECT 3.4650 0.9600 3.5650 1.1350 ;
        RECT 0.7250 0.6600 1.8000 0.7600 ;
        RECT 0.7250 0.7600 0.8150 1.2800 ;
    END
    ANTENNAGATEAREA 0.348 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 0.8500 1.6000 0.9500 ;
        RECT 1.0100 0.9500 1.1800 1.0200 ;
        RECT 1.5000 0.9500 1.6000 1.0500 ;
        RECT 1.0650 1.0200 1.1800 1.4800 ;
        RECT 1.5000 1.0500 1.8850 1.1100 ;
        RECT 0.4350 1.4800 1.7200 1.5700 ;
        RECT 1.5000 1.1100 2.6200 1.1400 ;
        RECT 1.6300 1.5700 1.7200 1.6950 ;
        RECT 0.4350 0.8400 0.5250 1.4800 ;
        RECT 1.5000 1.1400 2.4000 1.1500 ;
        RECT 2.3100 1.0500 2.6200 1.1100 ;
        RECT 1.6300 1.6950 2.7700 1.7850 ;
        RECT 1.7750 1.1500 2.4000 1.2100 ;
        RECT 2.6800 1.5700 2.7700 1.6950 ;
        RECT 2.6800 1.4800 3.3250 1.5700 ;
        RECT 3.2350 1.0500 3.3250 1.4800 ;
    END
    ANTENNAGATEAREA 0.348 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8100 1.4500 2.5900 1.5500 ;
        RECT 1.8100 1.3900 1.9000 1.4500 ;
        RECT 2.4900 1.3500 2.5900 1.4500 ;
        RECT 1.3100 1.3000 1.9000 1.3900 ;
        RECT 2.4900 1.2500 2.8400 1.3500 ;
        RECT 1.3100 1.0600 1.4000 1.3000 ;
        RECT 2.7350 1.1500 2.8400 1.2500 ;
        RECT 2.7350 1.0500 3.1050 1.1500 ;
    END
    ANTENNAGATEAREA 0.348 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 2.0800 1.8950 2.2500 2.0800 ;
        RECT 0.7350 1.8400 0.8350 2.0800 ;
        RECT 3.6350 1.8400 3.7350 2.0800 ;
        RECT 4.1550 1.8000 4.2550 2.0800 ;
        RECT 4.6700 1.8000 4.7800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.8900 0.6700 3.8000 0.7600 ;
      RECT 3.7100 0.7600 3.8000 1.6600 ;
      RECT 2.8600 1.6600 3.8000 1.7500 ;
      RECT 0.0800 0.7500 0.1700 1.6600 ;
      RECT 0.0800 0.6600 0.5400 0.7500 ;
      RECT 0.4500 0.5700 0.5400 0.6600 ;
      RECT 1.3600 1.7500 1.5300 1.9500 ;
      RECT 0.0800 1.6600 1.5300 1.7500 ;
      RECT 0.4500 0.4800 1.9800 0.5700 ;
      RECT 1.8900 0.5700 1.9800 0.6700 ;
      RECT 2.2950 0.4550 2.4650 0.6700 ;
      RECT 2.8150 0.4550 2.9850 0.6700 ;
      RECT 2.8600 1.7500 3.0300 1.9500 ;
      RECT 3.3350 0.4550 3.5050 0.6700 ;
  END
END OR3_X4M_A12TH

MACRO OR3_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.4200 0.3200 0.5200 0.5750 ;
        RECT 0.9400 0.3200 1.0400 0.5750 ;
        RECT 1.4600 0.3200 1.5600 0.5750 ;
        RECT 1.9800 0.3200 2.0800 0.5750 ;
        RECT 2.5000 0.3200 2.6000 0.5750 ;
        RECT 3.0200 0.3200 3.1200 0.5750 ;
        RECT 3.5400 0.3200 3.6400 0.5750 ;
        RECT 3.8200 0.3200 3.9200 0.5750 ;
        RECT 4.3400 0.3200 4.4400 0.5750 ;
        RECT 4.8600 0.3200 4.9600 0.5750 ;
        RECT 5.3800 0.3200 5.4800 0.5750 ;
        RECT 5.8500 0.3200 5.9500 0.5750 ;
        RECT 6.3700 0.3200 6.4700 0.6450 ;
        RECT 6.8900 0.3200 6.9900 0.6450 ;
        RECT 7.4100 0.3200 7.5100 0.6450 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 5.8500 1.7700 5.9500 2.0800 ;
        RECT 6.3700 1.7700 6.4700 2.0800 ;
        RECT 6.8900 1.7700 6.9900 2.0800 ;
        RECT 7.4100 1.7700 7.5100 2.0800 ;
        RECT 0.6800 1.7100 0.7800 2.0800 ;
        RECT 1.2000 1.7100 1.3000 2.0800 ;
        RECT 1.7200 1.7100 1.8200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 0.9400 7.3500 1.2700 ;
        RECT 6.1100 1.2700 7.3500 1.3700 ;
        RECT 6.1100 0.8400 7.3500 0.9400 ;
        RECT 6.1100 1.3700 6.2100 1.7300 ;
        RECT 6.6300 1.3700 6.7300 1.7200 ;
        RECT 7.1500 1.3700 7.2500 1.7200 ;
        RECT 6.1100 0.4900 6.2100 0.8400 ;
        RECT 6.6300 0.4900 6.7300 0.8400 ;
        RECT 7.1500 0.4900 7.2500 0.8400 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8500 1.6800 0.9500 ;
    END
    ANTENNAGATEAREA 0.5184 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4400 0.8500 3.2400 0.9500 ;
    END
    ANTENNAGATEAREA 0.5184 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2300 0.8500 5.0800 0.9500 ;
    END
    ANTENNAGATEAREA 0.5184 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4250 1.3000 3.6350 1.3900 ;
      RECT 1.9850 1.3900 2.0750 1.7000 ;
      RECT 2.5050 1.3900 2.5950 1.7000 ;
      RECT 3.0250 1.3900 3.1150 1.7000 ;
      RECT 3.5450 1.3900 3.6350 1.7000 ;
      RECT 0.4250 1.3900 0.5150 1.7200 ;
      RECT 0.9450 1.3900 1.0350 1.7150 ;
      RECT 1.4650 1.3900 1.5550 1.7150 ;
      RECT 2.2450 1.8300 5.4750 1.9200 ;
      RECT 2.2450 1.5100 2.3350 1.8300 ;
      RECT 2.7650 1.5100 2.8550 1.8300 ;
      RECT 3.2850 1.5100 3.3750 1.8300 ;
      RECT 3.8250 1.5100 3.9150 1.8300 ;
      RECT 4.3450 1.5100 4.4350 1.8300 ;
      RECT 4.8650 1.5100 4.9550 1.8300 ;
      RECT 5.3850 1.5100 5.4750 1.8300 ;
      RECT 5.8550 1.0600 6.9200 1.1500 ;
      RECT 4.6050 1.3900 4.6950 1.7000 ;
      RECT 4.6000 0.4600 4.7000 0.6650 ;
      RECT 5.1250 1.3900 5.2150 1.7000 ;
      RECT 5.1200 0.4600 5.2200 0.6650 ;
      RECT 4.0850 1.3000 5.9450 1.3900 ;
      RECT 5.8550 1.1500 5.9450 1.3000 ;
      RECT 5.8550 0.7550 5.9450 1.0600 ;
      RECT 0.6850 0.6650 5.9450 0.7550 ;
      RECT 2.7600 0.4600 2.8600 0.6650 ;
      RECT 3.2800 0.4600 3.3800 0.6650 ;
      RECT 4.0850 1.3900 4.1750 1.7000 ;
      RECT 4.0800 0.4600 4.1800 0.6650 ;
      RECT 1.2000 0.4600 1.3000 0.6650 ;
      RECT 1.7200 0.4600 1.8200 0.6650 ;
      RECT 2.2400 0.4600 2.3400 0.6650 ;
      RECT 0.6850 0.4600 0.7750 0.6650 ;
  END
END OR3_X6M_A12TH

MACRO OR3_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 9.8450 0.3200 ;
        RECT 0.4200 0.3200 0.5200 0.5700 ;
        RECT 0.9400 0.3200 1.0400 0.5700 ;
        RECT 1.4600 0.3200 1.5600 0.5700 ;
        RECT 1.9800 0.3200 2.0800 0.5700 ;
        RECT 2.5000 0.3200 2.6000 0.5700 ;
        RECT 2.7800 0.3200 2.8800 0.5700 ;
        RECT 3.3000 0.3200 3.4000 0.5700 ;
        RECT 3.8200 0.3200 3.9200 0.5700 ;
        RECT 4.3400 0.3200 4.4400 0.5700 ;
        RECT 4.8600 0.3200 4.9600 0.5700 ;
        RECT 5.3800 0.3200 5.4800 0.5700 ;
        RECT 5.9000 0.3200 6.0000 0.5700 ;
        RECT 6.4200 0.3200 6.5200 0.5700 ;
        RECT 6.9400 0.3200 7.0400 0.5700 ;
        RECT 7.5300 0.3200 7.6300 0.5800 ;
        RECT 8.0500 0.3200 8.1500 0.6450 ;
        RECT 8.5700 0.3200 8.6700 0.6450 ;
        RECT 9.0900 0.3200 9.1900 0.6450 ;
        RECT 9.6100 0.3200 9.7100 0.6450 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.8500 4.5000 0.9500 ;
    END
    ANTENNAGATEAREA 0.6984 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3000 0.8500 6.5000 0.9500 ;
    END
    ANTENNAGATEAREA 0.6984 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 9.8450 2.7200 ;
        RECT 0.4200 1.7700 0.5200 2.0800 ;
        RECT 0.9400 1.7700 1.0400 2.0800 ;
        RECT 1.4600 1.7700 1.5600 2.0800 ;
        RECT 1.9800 1.7700 2.0800 2.0800 ;
        RECT 2.5000 1.7700 2.6000 2.0800 ;
        RECT 7.5300 1.7700 7.6300 2.0800 ;
        RECT 8.0500 1.7700 8.1500 2.0800 ;
        RECT 8.5700 1.7700 8.6700 2.0800 ;
        RECT 9.0900 1.7700 9.1900 2.0800 ;
        RECT 9.6100 1.7700 9.7100 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 0.8500 2.1000 0.9500 ;
    END
    ANTENNAGATEAREA 0.6984 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.8250 1.3850 8.9650 1.7200 ;
        RECT 7.7750 1.2550 9.5600 1.3850 ;
        RECT 7.7750 1.3850 7.9050 1.7300 ;
        RECT 8.2950 1.3850 8.4250 1.7200 ;
        RECT 9.3350 1.3850 9.4650 1.7200 ;
        RECT 9.4300 0.9550 9.5600 1.2550 ;
        RECT 7.7750 0.8250 9.5600 0.9550 ;
        RECT 7.7750 0.4900 7.9050 0.8250 ;
        RECT 8.2950 0.4900 8.4250 0.8250 ;
        RECT 8.8150 0.4900 8.9450 0.8250 ;
        RECT 9.3350 0.4900 9.4650 0.8250 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 7.4550 1.0600 9.1000 1.1500 ;
      RECT 5.6450 1.3900 5.7350 1.7000 ;
      RECT 5.6400 0.4650 5.7400 0.6700 ;
      RECT 6.1650 1.3900 6.2550 1.7000 ;
      RECT 6.1600 0.4650 6.2600 0.6700 ;
      RECT 6.6850 1.3900 6.7750 1.7000 ;
      RECT 6.6800 0.4650 6.7800 0.6700 ;
      RECT 5.1250 1.3000 7.5550 1.3900 ;
      RECT 7.4650 1.1500 7.5550 1.3000 ;
      RECT 7.4650 0.7600 7.5550 1.0600 ;
      RECT 0.6850 0.6700 7.5550 0.7600 ;
      RECT 3.5600 0.4650 3.6600 0.6700 ;
      RECT 4.0800 0.4650 4.1800 0.6700 ;
      RECT 4.6000 0.4650 4.7000 0.6700 ;
      RECT 5.1250 1.3900 5.2150 1.7000 ;
      RECT 5.1200 0.4650 5.2200 0.6700 ;
      RECT 1.2000 0.4650 1.3000 0.6700 ;
      RECT 1.7200 0.4650 1.8200 0.6700 ;
      RECT 2.2400 0.4650 2.3400 0.6700 ;
      RECT 3.0400 0.4650 3.1400 0.6700 ;
      RECT 0.6850 0.4650 0.7750 0.6700 ;
      RECT 0.6850 1.3900 0.7750 1.7200 ;
      RECT 0.6850 1.3000 4.6950 1.3900 ;
      RECT 1.2050 1.3900 1.2950 1.7150 ;
      RECT 1.7250 1.3900 1.8150 1.7150 ;
      RECT 2.2450 1.3900 2.3350 1.7000 ;
      RECT 3.0450 1.3900 3.1350 1.7000 ;
      RECT 3.5650 1.3900 3.6550 1.7000 ;
      RECT 4.0850 1.3900 4.1750 1.7000 ;
      RECT 4.6050 1.3900 4.6950 1.7000 ;
      RECT 2.7850 1.8300 7.0350 1.9200 ;
      RECT 2.7850 1.5100 2.8750 1.8300 ;
      RECT 3.3050 1.5100 3.3950 1.8300 ;
      RECT 3.8250 1.5100 3.9150 1.8300 ;
      RECT 4.3450 1.5100 4.4350 1.8300 ;
      RECT 4.8650 1.5100 4.9550 1.8300 ;
      RECT 5.3850 1.5100 5.4750 1.8300 ;
      RECT 5.9050 1.5100 5.9950 1.8300 ;
      RECT 6.4250 1.5100 6.5150 1.8300 ;
      RECT 6.9450 1.5100 7.0350 1.8300 ;
  END
END OR3_X8M_A12TH

MACRO OR4_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6900 ;
        RECT 0.5950 0.3200 0.6950 0.6950 ;
        RECT 1.2900 0.3200 1.3900 0.7650 ;
        RECT 1.8250 0.3200 1.9250 0.7650 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7800 0.1650 0.9400 ;
        RECT 0.0500 0.9400 0.2750 1.1500 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0100 0.5500 1.2350 ;
        RECT 0.3050 1.2350 0.5500 1.3350 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8400 1.0900 1.9500 1.5900 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1850 1.4500 1.5100 1.5500 ;
        RECT 1.4200 1.5500 1.5100 1.6000 ;
        RECT 1.4200 1.3900 1.5100 1.4500 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8450 0.8500 1.1900 0.9500 ;
        RECT 1.0050 0.9500 1.0950 1.6950 ;
        RECT 0.8450 0.5800 0.9350 0.8500 ;
        RECT 1.0050 1.6950 1.1250 1.9050 ;
    END
    ANTENNADIFFAREA 0.1236 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.7700 1.8700 0.8700 2.0800 ;
        RECT 1.3500 1.6900 1.4500 2.0800 ;
        RECT 0.0750 1.4100 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2850 0.5600 0.4900 0.6600 ;
      RECT 0.4000 0.6600 0.4900 0.8050 ;
      RECT 0.4000 0.8050 0.7450 0.8950 ;
      RECT 0.5700 1.5250 0.6700 1.8000 ;
      RECT 0.5700 1.4300 0.7450 1.5250 ;
      RECT 0.6550 1.2850 0.7450 1.4300 ;
      RECT 0.6550 0.8950 0.7450 1.0750 ;
      RECT 0.6550 1.0750 0.9150 1.2850 ;
      RECT 1.7750 1.7900 1.9450 1.9900 ;
      RECT 1.6200 1.7000 1.9450 1.7900 ;
      RECT 1.1900 1.0700 1.2800 1.1900 ;
      RECT 1.6200 1.2800 1.7100 1.7000 ;
      RECT 1.1900 1.1900 1.7100 1.2800 ;
      RECT 1.6200 0.7650 1.7100 1.1900 ;
      RECT 1.5700 0.6750 1.7100 0.7650 ;
      RECT 1.5700 0.5550 1.6600 0.6750 ;
  END
END OR4_X0P5M_A12TH

MACRO OR4_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.5800 0.3200 0.6700 0.8650 ;
        RECT 0.0800 0.3200 0.1700 0.9850 ;
        RECT 1.2750 0.3200 1.3750 0.7200 ;
        RECT 1.8250 0.3200 1.9250 0.7350 ;
        RECT 0.5800 0.8650 0.7700 0.9550 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7800 0.6500 1.1050 0.7500 ;
        RECT 1.0150 0.7500 1.1050 1.6000 ;
        RECT 0.7800 0.4200 0.9500 0.6500 ;
        RECT 1.0150 1.6000 1.1700 1.6900 ;
        RECT 1.0800 1.6900 1.1700 1.9900 ;
    END
    ANTENNADIFFAREA 0.1752 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4500 0.3900 1.5800 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1700 1.2500 0.5900 1.3500 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8100 1.3500 1.0500 ;
        RECT 1.2500 1.0500 1.5500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0150 1.9500 1.2500 ;
        RECT 1.8400 0.8450 1.9500 1.0150 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.7800 1.7800 0.9500 2.0800 ;
        RECT 0.0900 1.7200 0.1800 2.0800 ;
        RECT 1.3400 1.6550 1.4300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.7850 0.4300 1.0500 ;
      RECT 0.3400 1.0500 0.7700 1.1400 ;
      RECT 0.5000 1.6000 0.7700 1.6900 ;
      RECT 0.5000 1.6900 0.6700 1.9850 ;
      RECT 0.6800 1.4500 0.7700 1.6000 ;
      RECT 0.6800 1.1400 0.7700 1.2400 ;
      RECT 0.6800 1.2400 0.9250 1.4500 ;
      RECT 1.8050 1.4850 1.8950 1.9900 ;
      RECT 1.2050 1.3950 1.8950 1.4850 ;
      RECT 1.6400 0.8600 1.7300 1.3950 ;
      RECT 1.5700 0.7700 1.7300 0.8600 ;
      RECT 1.5700 0.5600 1.6600 0.7700 ;
      RECT 1.2050 1.2600 1.2950 1.3950 ;
  END
END OR4_X0P7M_A12TH

MACRO OR4_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5450 ;
        RECT 0.5950 0.3200 0.6950 0.5400 ;
        RECT 1.2900 0.3200 1.3900 0.5900 ;
        RECT 1.8250 0.3200 1.9250 0.9100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.3250 1.8800 1.4350 2.0800 ;
        RECT 0.7850 1.7350 0.8850 2.0800 ;
        RECT 0.0750 1.5550 0.1750 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.2350 1.7600 1.5050 ;
        RECT 1.6500 1.0650 1.8150 1.2350 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0550 1.5600 1.5050 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8300 0.8700 1.1450 0.9900 ;
        RECT 1.0500 0.9900 1.1450 1.8350 ;
        RECT 0.8300 0.7900 0.9500 0.8700 ;
    END
    ANTENNADIFFAREA 0.238625 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8950 0.1600 1.3050 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9900 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.6450 1.0950 0.9450 1.2150 ;
      RECT 0.5350 1.5700 0.6350 1.8900 ;
      RECT 0.5350 1.4800 0.7350 1.5700 ;
      RECT 0.6450 1.2150 0.7350 1.4800 ;
      RECT 0.6450 0.7200 0.7350 1.0950 ;
      RECT 0.3400 0.6300 0.7350 0.7200 ;
      RECT 0.3400 0.4400 0.4300 0.6300 ;
      RECT 1.8300 1.7700 1.9200 1.8850 ;
      RECT 1.2350 1.6800 1.9200 1.7700 ;
      RECT 1.2350 0.8200 1.7150 0.9100 ;
      RECT 1.2350 0.9100 1.3250 1.6800 ;
  END
END OR4_X1M_A12TH

MACRO OR4_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.4850 ;
        RECT 0.5400 0.3200 0.7500 0.3850 ;
        RECT 1.4500 0.3200 1.6600 0.3850 ;
        RECT 2.0250 0.3200 2.1250 0.5650 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8100 1.7550 1.2300 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.5150 1.8250 1.6250 2.0800 ;
        RECT 0.9850 1.8150 1.0850 2.0800 ;
        RECT 0.5350 1.7900 0.6350 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0250 0.8850 2.1500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8350 0.1600 1.3050 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9900 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.4450 1.1500 0.7400 ;
        RECT 0.8550 0.7400 1.1500 0.8400 ;
        RECT 0.8550 0.8400 0.9550 1.2500 ;
        RECT 0.8550 1.2500 1.3450 1.3500 ;
        RECT 1.2450 1.3500 1.3450 1.4800 ;
    END
    ANTENNADIFFAREA 0.285 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5900 1.5250 1.6800 ;
      RECT 1.4350 1.0450 1.5250 1.5900 ;
      RECT 0.0750 1.6800 0.1750 1.9800 ;
      RECT 0.6750 0.5700 0.7650 1.5900 ;
      RECT 0.2750 0.4800 0.7650 0.5700 ;
      RECT 2.0300 1.6750 2.1200 1.9750 ;
      RECT 1.8450 1.5850 2.1200 1.6750 ;
      RECT 1.8450 0.5700 1.9350 1.5850 ;
      RECT 1.2550 0.4800 1.9350 0.5700 ;
      RECT 1.2550 0.5700 1.3450 1.0050 ;
      RECT 1.0750 1.0050 1.3450 1.0950 ;
  END
END OR4_X1P4M_A12TH

MACRO OR4_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5700 ;
        RECT 0.5950 0.3200 0.6950 0.5550 ;
        RECT 1.8250 0.3200 1.9250 0.5850 ;
        RECT 2.4850 0.3200 2.5850 0.4250 ;
        RECT 3.0250 0.3200 3.1250 0.5600 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1350 1.0400 2.9650 1.1500 ;
        RECT 2.8750 1.1500 2.9650 1.2100 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3800 0.8500 2.8000 0.9500 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.1500 1.7500 1.5200 ;
        RECT 1.3050 1.5200 1.9250 1.6200 ;
        RECT 1.3400 1.0500 1.7500 1.1500 ;
        RECT 1.3050 1.6200 1.4050 1.9550 ;
        RECT 1.8250 1.6200 1.9250 1.9550 ;
        RECT 1.3400 0.9550 1.4400 1.0500 ;
        RECT 1.2700 0.6650 1.4400 0.9550 ;
    END
    ANTENNADIFFAREA 0.402 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.0500 1.0950 1.1500 ;
        RECT 0.2350 0.9400 0.3350 1.0500 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 0.8500 0.8800 0.9600 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.5650 1.7100 1.6650 2.0800 ;
        RECT 0.0750 1.5600 0.1750 2.0800 ;
        RECT 1.0450 1.5600 1.1450 2.0800 ;
        RECT 2.0850 1.5600 2.1850 2.0800 ;
        RECT 3.0250 1.5600 3.1250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.3000 1.4600 1.3900 ;
      RECT 1.2500 1.2600 1.4600 1.3000 ;
      RECT 0.5950 1.3900 0.6950 1.8850 ;
      RECT 0.0550 0.6700 0.4300 0.7600 ;
      RECT 0.3400 0.4800 0.4300 0.6700 ;
      RECT 0.0550 0.7600 0.1450 1.3000 ;
      RECT 1.5700 0.8200 2.1800 0.9100 ;
      RECT 2.0900 0.4800 2.1800 0.8200 ;
      RECT 1.0500 0.4800 1.6600 0.5700 ;
      RECT 1.5700 0.5700 1.6600 0.8200 ;
      RECT 1.0500 0.5700 1.1400 0.9100 ;
      RECT 1.8650 1.3200 3.1550 1.4100 ;
      RECT 3.0650 0.7600 3.1550 1.3200 ;
      RECT 2.7700 0.6700 3.1550 0.7600 ;
      RECT 1.8650 1.2550 2.0450 1.3200 ;
      RECT 2.5350 1.4100 2.6350 1.8850 ;
      RECT 2.7700 0.4700 2.8600 0.6700 ;
  END
END OR4_X2M_A12TH

MACRO OR4_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.5650 ;
        RECT 0.6100 0.3200 0.7100 0.5650 ;
        RECT 2.1100 0.3200 2.2100 0.6300 ;
        RECT 2.6300 0.3200 2.7300 0.6300 ;
        RECT 3.0900 0.3200 3.1900 0.6300 ;
        RECT 3.6100 0.3200 3.7100 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 1.5900 1.8150 1.6900 2.0800 ;
        RECT 2.1100 1.8150 2.2100 2.0800 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 1.0700 1.7700 1.1700 2.0800 ;
        RECT 2.6300 1.7700 2.7300 2.0800 ;
        RECT 3.6100 1.7700 3.7100 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 1.1200 1.3500 ;
        RECT 0.2500 0.9700 0.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1500 1.9500 1.6200 ;
        RECT 1.3300 1.6200 2.4700 1.7200 ;
        RECT 1.6300 1.0500 1.9500 1.1500 ;
        RECT 1.3300 1.7200 1.4300 1.9900 ;
        RECT 1.8550 1.7200 1.9450 1.9900 ;
        RECT 2.3700 1.7200 2.4700 1.9900 ;
        RECT 1.6300 0.9800 1.7300 1.0500 ;
        RECT 1.0750 0.8900 1.7300 0.9800 ;
        RECT 1.5550 0.6650 1.7300 0.8900 ;
        RECT 1.0750 0.5600 1.1650 0.8900 ;
    END
    ANTENNADIFFAREA 0.66075 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8950 1.0500 3.3450 1.1500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.9800 3.5500 1.2600 ;
        RECT 2.7000 1.2600 3.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END D
  OBS
    LAYER M1 ;
      RECT 2.0800 1.4400 3.7500 1.5300 ;
      RECT 3.6600 0.8550 3.7500 1.4400 ;
      RECT 3.3550 0.7650 3.7500 0.8550 ;
      RECT 2.0800 1.3950 2.4900 1.4400 ;
      RECT 3.0900 1.5300 3.1900 1.8700 ;
      RECT 3.3550 0.4850 3.4450 0.7650 ;
      RECT 0.0500 1.4400 1.7200 1.5300 ;
      RECT 1.3100 1.3950 1.7200 1.4400 ;
      RECT 0.6100 1.5300 0.7100 1.8700 ;
      RECT 0.0500 0.6900 0.4450 0.7800 ;
      RECT 0.3550 0.4100 0.4450 0.6900 ;
      RECT 0.0500 0.7800 0.1400 1.4400 ;
      RECT 1.8550 0.8150 2.4650 0.9050 ;
      RECT 2.3750 0.4700 2.4650 0.8150 ;
      RECT 1.8550 0.5700 1.9450 0.8150 ;
      RECT 1.2750 0.4800 1.9450 0.5700 ;
  END
END OR4_X3M_A12TH

MACRO OR4_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.4950 0.3200 0.6000 0.5700 ;
        RECT 1.0300 0.3200 1.1300 0.5600 ;
        RECT 1.5750 0.3200 1.6750 0.5450 ;
        RECT 2.5550 0.3200 2.6550 0.5450 ;
        RECT 3.6350 0.3200 3.7350 0.5450 ;
        RECT 4.2900 0.3200 4.3900 0.5450 ;
        RECT 4.8100 0.3200 4.9100 0.5450 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.0500 1.2750 1.1500 ;
        RECT 0.2350 1.1500 0.3250 1.3100 ;
    END
    ANTENNAGATEAREA 0.1776 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.9500 3.7500 1.2700 ;
        RECT 3.5350 1.2700 3.7500 1.3600 ;
        RECT 3.6500 0.8500 4.4350 0.9500 ;
    END
    ANTENNAGATEAREA 0.1767 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.2500 1.4850 1.3500 ;
        RECT 1.3850 1.1450 1.4850 1.2500 ;
    END
    ANTENNAGATEAREA 0.1776 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7300 1.6500 3.1850 1.7500 ;
        RECT 1.7300 1.7500 1.9000 1.9550 ;
        RECT 2.2600 1.7500 2.4300 1.9550 ;
        RECT 2.7800 1.7500 2.9500 1.9550 ;
        RECT 3.0950 0.9250 3.1850 1.6500 ;
        RECT 1.9750 0.8250 3.1850 0.9250 ;
    END
    ANTENNADIFFAREA 0.8143 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2400 1.2000 4.3500 1.4500 ;
        RECT 3.2750 1.4500 4.3500 1.5500 ;
        RECT 4.2400 1.1900 4.7350 1.2000 ;
        RECT 3.2750 1.2450 3.3650 1.4500 ;
        RECT 3.9000 1.1000 4.7350 1.1900 ;
        RECT 4.6450 0.8300 4.7350 1.1000 ;
    END
    ANTENNAGATEAREA 0.1767 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 2.0350 1.8400 2.1350 2.0800 ;
        RECT 2.5550 1.8400 2.6550 2.0800 ;
        RECT 3.1150 1.8400 3.2150 2.0800 ;
        RECT 4.0750 1.8400 4.1750 2.0800 ;
        RECT 0.5700 1.8000 0.6700 2.0800 ;
        RECT 1.4950 1.8000 1.5950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.4400 3.0050 1.5300 ;
      RECT 2.9150 1.0700 3.0050 1.4400 ;
      RECT 0.0500 1.5300 0.1700 1.9100 ;
      RECT 0.0500 0.7600 0.1400 1.4400 ;
      RECT 0.7600 0.4450 0.8600 0.6700 ;
      RECT 0.0500 0.6700 1.3900 0.7600 ;
      RECT 1.2900 0.4450 1.3900 0.6700 ;
      RECT 1.0300 1.5300 1.1300 1.9150 ;
      RECT 2.0050 1.2000 2.1750 1.4400 ;
      RECT 3.5700 1.6400 4.9350 1.7300 ;
      RECT 4.8450 0.7300 4.9350 1.6400 ;
      RECT 3.4250 0.7250 4.9350 0.7300 ;
      RECT 1.6850 0.6400 4.9350 0.7250 ;
      RECT 1.6850 0.7250 1.7750 1.0200 ;
      RECT 1.6850 1.1100 1.7800 1.2650 ;
      RECT 1.6850 1.0200 2.7900 1.1100 ;
      RECT 2.4200 1.1100 2.7900 1.1800 ;
      RECT 3.4250 0.7300 3.5150 1.0350 ;
      RECT 3.3200 1.0350 3.5150 1.1350 ;
      RECT 1.6850 0.6350 4.1650 0.6400 ;
      RECT 3.9950 0.4850 4.1650 0.6350 ;
      RECT 3.5700 1.7300 3.7400 1.9550 ;
      RECT 4.5250 1.7300 4.6950 1.9550 ;
      RECT 4.5150 0.4850 4.6850 0.6400 ;
  END
END OR4_X4M_A12TH

MACRO OR4_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.8950 0.3200 0.9950 0.5450 ;
        RECT 1.4350 0.3200 1.5400 0.6000 ;
        RECT 1.9700 0.3200 2.1400 0.5200 ;
        RECT 3.0550 0.3200 3.1550 0.5450 ;
        RECT 4.0950 0.3200 4.1950 0.5450 ;
        RECT 5.1350 0.3200 5.2350 0.6150 ;
        RECT 5.5850 0.3200 5.6850 0.6200 ;
        RECT 6.1050 0.3200 6.2050 0.6200 ;
        RECT 6.6250 0.3200 6.7250 0.6200 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 0.8500 0.9900 0.9650 ;
        RECT 0.4000 0.9650 1.9400 1.0750 ;
    END
    ANTENNAGATEAREA 0.2616 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4100 1.0500 6.3750 1.1500 ;
        RECT 5.4100 1.1500 5.5100 1.2700 ;
        RECT 5.1650 1.2700 5.5100 1.3600 ;
    END
    ANTENNAGATEAREA 0.2616 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.2500 1.6950 1.3500 ;
    END
    ANTENNAGATEAREA 0.2616 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2750 1.6200 4.7750 1.7500 ;
        RECT 2.2750 1.7500 2.3750 1.9900 ;
        RECT 2.7950 1.7500 2.8950 1.9900 ;
        RECT 3.3150 1.7500 3.4150 1.9900 ;
        RECT 3.8350 1.7500 3.9350 1.9900 ;
        RECT 4.3550 1.7500 4.4550 1.9900 ;
        RECT 4.6850 0.9550 4.7750 1.6200 ;
        RECT 4.2450 0.8650 4.7750 0.9550 ;
        RECT 4.2450 0.9550 4.3350 1.2600 ;
        RECT 3.7550 1.2600 4.3350 1.3500 ;
        RECT 3.7550 0.9600 3.8450 1.2600 ;
        RECT 3.2650 0.8600 3.8450 0.9600 ;
        RECT 3.2650 0.9600 3.3550 1.2600 ;
        RECT 2.8050 1.2600 3.3550 1.3500 ;
        RECT 2.8050 0.9600 2.8950 1.2600 ;
        RECT 2.4800 0.8650 2.8950 0.9600 ;
    END
    ANTENNADIFFAREA 1.25295 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6600 1.2500 6.5750 1.3500 ;
        RECT 5.6600 1.3500 5.7500 1.4500 ;
        RECT 6.4850 1.1400 6.5750 1.2500 ;
        RECT 4.8650 1.4500 5.7500 1.5400 ;
        RECT 4.8650 1.2100 4.9550 1.4500 ;
    END
    ANTENNAGATEAREA 0.2616 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 2.5000 1.8650 2.6700 2.0800 ;
        RECT 3.0200 1.8650 3.1900 2.0800 ;
        RECT 3.5400 1.8650 3.7100 2.0800 ;
        RECT 4.0600 1.8650 4.2300 2.0800 ;
        RECT 4.6450 1.8650 4.8150 2.0800 ;
        RECT 5.6850 1.8400 5.7850 2.0800 ;
        RECT 6.6250 1.8300 6.7250 2.0800 ;
        RECT 0.0750 1.8100 0.1750 2.0800 ;
        RECT 0.9950 1.8100 1.0950 2.0800 ;
        RECT 1.9900 1.8100 2.0900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.6250 1.4400 4.5150 1.5300 ;
      RECT 4.4250 1.2100 4.5150 1.4400 ;
      RECT 4.4250 1.1200 4.5950 1.2100 ;
      RECT 0.1900 0.7450 0.2800 1.4600 ;
      RECT 0.5350 1.5500 0.6350 1.8650 ;
      RECT 0.1900 0.6550 1.2500 0.7450 ;
      RECT 1.1600 0.7450 1.2500 0.7650 ;
      RECT 1.1600 0.4850 1.2500 0.6550 ;
      RECT 1.5000 1.5500 1.6000 1.8650 ;
      RECT 1.1600 0.7650 1.7950 0.8550 ;
      RECT 1.6950 0.4850 1.7950 0.7650 ;
      RECT 0.1900 1.4600 2.0750 1.5500 ;
      RECT 1.9850 1.3700 2.0750 1.4600 ;
      RECT 1.9850 1.2800 2.7150 1.3700 ;
      RECT 2.6250 1.3700 2.7150 1.4400 ;
      RECT 3.4450 1.3000 3.5350 1.4400 ;
      RECT 3.4450 1.2100 3.6450 1.3000 ;
      RECT 5.1900 1.6300 6.7550 1.7200 ;
      RECT 6.6650 0.8700 6.7550 1.6300 ;
      RECT 4.9350 0.7800 6.7550 0.8700 ;
      RECT 2.3000 0.7250 2.3900 1.0800 ;
      RECT 2.0350 1.0800 2.3900 1.1700 ;
      RECT 3.0850 0.7250 3.1750 1.0800 ;
      RECT 3.0050 1.0800 3.1750 1.1700 ;
      RECT 4.0450 0.7250 4.1350 1.0800 ;
      RECT 3.9550 1.0800 4.1350 1.1700 ;
      RECT 4.9350 0.7250 5.0250 0.7800 ;
      RECT 2.3000 0.6350 5.0250 0.7250 ;
      RECT 5.1900 1.7200 5.3600 1.9200 ;
      RECT 5.0850 0.8700 5.1750 1.1800 ;
      RECT 5.8450 0.4600 5.9450 0.7800 ;
      RECT 6.1100 1.7200 6.2800 1.9550 ;
      RECT 6.3650 0.4600 6.4600 0.7800 ;
  END
END OR4_X6M_A12TH

MACRO OR4_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 9.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5600 ;
        RECT 0.5950 0.3200 0.6950 0.5350 ;
        RECT 1.1150 0.3200 1.2150 0.5350 ;
        RECT 1.6350 0.3200 1.7350 0.5350 ;
        RECT 2.1550 0.3200 2.2550 0.5350 ;
        RECT 2.6500 0.3200 2.8200 0.4550 ;
        RECT 3.6000 0.3200 3.7050 0.5450 ;
        RECT 4.6250 0.3200 4.7250 0.5450 ;
        RECT 5.6650 0.3200 5.7650 0.5450 ;
        RECT 6.5650 0.3200 6.7400 0.4700 ;
        RECT 7.1450 0.3200 7.2450 0.5350 ;
        RECT 7.6650 0.3200 7.7650 0.5350 ;
        RECT 8.1850 0.3200 8.2850 0.5350 ;
        RECT 8.7050 0.3200 8.8050 0.5350 ;
        RECT 9.2250 0.3200 9.3250 0.5450 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2650 0.8500 2.3750 0.9500 ;
        RECT 0.2650 0.9500 0.3550 1.1200 ;
    END
    ANTENNAGATEAREA 0.3555 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.8500 8.9350 0.9500 ;
        RECT 6.8150 0.9500 6.9050 1.0400 ;
    END
    ANTENNAGATEAREA 0.3555 ;
  END D

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0500 2.5250 1.1550 ;
        RECT 2.4350 1.1550 2.5250 1.2550 ;
    END
    ANTENNAGATEAREA 0.3555 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4350 1.7500 6.5650 1.9900 ;
        RECT 2.8050 1.6200 6.5650 1.7500 ;
        RECT 2.8050 1.7500 2.9050 1.9900 ;
        RECT 3.3250 1.7500 3.4250 1.9900 ;
        RECT 3.8450 1.7500 3.9450 1.9900 ;
        RECT 4.3650 1.7500 4.4650 1.9900 ;
        RECT 4.8850 1.7500 4.9850 1.9900 ;
        RECT 5.4000 1.7500 5.5050 1.9900 ;
        RECT 5.9200 1.7500 6.0250 1.9900 ;
        RECT 6.3550 1.6100 6.5650 1.6200 ;
        RECT 6.3550 0.9900 6.4850 1.6100 ;
        RECT 5.9100 0.8600 6.4850 0.9900 ;
        RECT 5.9100 0.9900 6.0400 1.2300 ;
        RECT 5.3900 1.2300 6.0400 1.3500 ;
        RECT 5.3900 0.9900 5.5200 1.2300 ;
        RECT 4.8800 0.8600 5.5200 0.9900 ;
        RECT 4.8800 0.9900 5.0100 1.2300 ;
        RECT 4.3600 1.2300 5.0100 1.3500 ;
        RECT 4.3600 0.9900 4.4900 1.2300 ;
        RECT 3.8900 0.8600 4.4900 0.9900 ;
        RECT 3.8900 0.9900 4.0200 1.2350 ;
        RECT 3.2350 1.2350 4.0200 1.3500 ;
        RECT 3.2350 0.9850 3.3650 1.2350 ;
        RECT 3.1100 0.8550 3.3650 0.9850 ;
    END
    ANTENNADIFFAREA 1.608 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0450 1.0500 9.1650 1.1500 ;
        RECT 9.0750 1.1500 9.1650 1.2550 ;
    END
    ANTENNAGATEAREA 0.3555 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 9.4450 2.7200 ;
        RECT 1.6150 2.0750 2.6400 2.0800 ;
        RECT 3.0300 1.8600 3.2000 2.0800 ;
        RECT 3.5500 1.8600 3.7200 2.0800 ;
        RECT 4.0700 1.8600 4.2400 2.0800 ;
        RECT 4.5900 1.8600 4.7600 2.0800 ;
        RECT 5.1100 1.8600 5.2800 2.0800 ;
        RECT 5.6300 1.8600 5.8000 2.0800 ;
        RECT 6.1500 1.8600 6.3200 2.0800 ;
        RECT 0.5950 1.7850 0.6950 2.0800 ;
        RECT 7.6650 1.7700 7.7600 2.0800 ;
        RECT 6.7000 1.7650 6.8050 2.0800 ;
        RECT 8.7050 1.7650 8.8050 2.0800 ;
        RECT 1.6150 1.7850 1.7150 2.0750 ;
        RECT 2.5400 1.7800 2.6400 2.0750 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.0800 1.4400 6.2450 1.5300 ;
      RECT 6.1550 1.2500 6.2450 1.4400 ;
      RECT 0.3350 0.4900 0.4350 0.6700 ;
      RECT 0.0800 0.7600 0.1700 1.4100 ;
      RECT 0.0800 1.5000 0.1750 1.8300 ;
      RECT 0.8550 0.4900 0.9550 0.6700 ;
      RECT 1.3750 0.4900 1.4750 0.6700 ;
      RECT 0.0800 1.4100 1.2150 1.5000 ;
      RECT 1.1150 1.5000 1.2150 1.8300 ;
      RECT 1.8950 0.4900 1.9950 0.6700 ;
      RECT 2.6150 0.7600 2.7050 1.4400 ;
      RECT 0.0800 0.6700 2.7050 0.7600 ;
      RECT 2.4150 0.6650 2.7050 0.6700 ;
      RECT 2.9550 1.3750 3.1250 1.4400 ;
      RECT 2.4150 0.4900 2.5150 0.6650 ;
      RECT 2.0800 1.5300 2.1750 1.8500 ;
      RECT 4.1300 1.2650 4.2300 1.4400 ;
      RECT 5.1200 1.2600 5.2200 1.4400 ;
      RECT 2.7950 0.6350 9.3450 0.7250 ;
      RECT 9.2550 0.7250 9.3450 1.4200 ;
      RECT 9.2300 1.4200 9.3450 1.7900 ;
      RECT 2.7950 0.7250 2.8850 1.2550 ;
      RECT 3.6700 0.7250 3.7600 1.0550 ;
      RECT 3.5250 1.0550 3.7600 1.1450 ;
      RECT 4.6800 0.7250 4.7700 1.0400 ;
      RECT 4.6000 1.0400 4.7700 1.1400 ;
      RECT 6.6050 0.7250 6.6950 1.3900 ;
      RECT 5.7100 0.7250 5.8000 1.0400 ;
      RECT 5.6300 1.0400 5.8000 1.1400 ;
      RECT 6.8850 0.4800 6.9850 0.6350 ;
      RECT 7.2050 1.4800 7.3050 1.8500 ;
      RECT 7.4050 0.4800 7.5050 0.6350 ;
      RECT 7.9250 0.4800 8.0250 0.6350 ;
      RECT 6.6050 1.3900 8.2850 1.4800 ;
      RECT 8.1850 1.4800 8.2850 1.8500 ;
      RECT 8.4450 0.4800 8.5450 0.6350 ;
      RECT 8.9650 0.4800 9.0650 0.6350 ;
  END
END OR4_X8M_A12TH

MACRO OR6_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5200 ;
        RECT 0.5600 0.3200 0.7300 0.4500 ;
        RECT 1.5350 0.3200 1.7050 0.9800 ;
        RECT 2.1100 0.3200 2.3200 0.7800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0550 1.0500 1.4450 1.1500 ;
        RECT 1.3450 1.1500 1.4450 1.5500 ;
        RECT 1.0550 0.7150 1.1450 1.0500 ;
        RECT 1.3450 1.5500 1.4650 1.7600 ;
    END
    ANTENNADIFFAREA 0.1313 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7700 0.1650 1.1900 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.7450 0.5500 1.1650 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9700 0.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END A

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5550 1.4500 1.8700 1.5500 ;
        RECT 1.7700 1.2600 1.8700 1.4500 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END F

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.4000 2.1500 1.6600 ;
        RECT 1.9950 1.1900 2.1500 1.4000 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END E

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.0700 2.3500 1.4950 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 1.6400 1.8550 1.8100 2.0800 ;
        RECT 0.1100 1.7000 0.2000 2.0800 ;
        RECT 1.1150 1.6500 1.2050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8550 1.3600 1.2500 1.4500 ;
      RECT 1.1600 1.2600 1.2500 1.3600 ;
      RECT 0.7500 1.6300 0.8400 1.9600 ;
      RECT 0.7500 1.5300 0.9450 1.6300 ;
      RECT 0.8550 1.4500 0.9450 1.5300 ;
      RECT 0.8550 0.6300 0.9450 1.3600 ;
      RECT 0.3600 0.6250 0.9450 0.6300 ;
      RECT 0.3600 0.5400 0.9900 0.6250 ;
      RECT 0.8200 0.4100 0.9900 0.5400 ;
      RECT 0.3600 0.5000 0.4700 0.5400 ;
      RECT 0.2800 0.4100 0.4700 0.5000 ;
      RECT 2.3500 1.7900 2.4400 1.9100 ;
      RECT 2.3500 1.7000 2.5400 1.7900 ;
      RECT 2.4500 0.9600 2.5400 1.7000 ;
      RECT 1.8100 0.8700 2.5400 0.9600 ;
      RECT 2.4300 0.6600 2.5400 0.8700 ;
      RECT 1.8100 0.9600 1.9000 1.0700 ;
      RECT 1.5350 1.0700 1.9000 1.1600 ;
      RECT 1.9100 0.6550 2.0000 0.8700 ;
      RECT 1.5350 1.1600 1.6250 1.3400 ;
  END
END OR6_X0P5M_A12TH

MACRO OR6_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.5400 0.3200 0.6300 0.5850 ;
        RECT 0.0800 0.3200 0.1700 0.7200 ;
        RECT 1.5200 0.3200 1.6900 0.5300 ;
        RECT 2.1550 0.3200 2.2450 0.5350 ;
        RECT 0.5400 0.5850 0.7500 0.6750 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.5250 ;
        RECT 1.2500 1.5250 1.4500 1.6150 ;
        RECT 1.0700 0.6000 1.3500 0.7000 ;
        RECT 1.3500 1.6150 1.4500 1.9550 ;
        RECT 1.0700 0.4100 1.2400 0.6000 ;
    END
    ANTENNADIFFAREA 0.1752 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9000 0.1600 1.3200 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.9950 0.5500 1.4150 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9950 0.7800 1.3550 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END A

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.1050 1.7600 1.5700 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END F

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7050 0.8500 2.1500 0.9500 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END E

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9700 2.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.1500 1.8200 0.2400 2.0800 ;
        RECT 1.6550 1.8200 1.7450 2.0800 ;
        RECT 1.0550 1.7050 1.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7900 1.5000 1.1500 1.5900 ;
      RECT 1.0600 0.8850 1.1500 1.5000 ;
      RECT 0.3400 0.7950 1.1500 0.8850 ;
      RECT 0.8600 0.7900 1.1500 0.7950 ;
      RECT 0.7900 1.5900 0.8800 1.9100 ;
      RECT 0.8600 0.5450 0.9500 0.7900 ;
      RECT 0.3400 0.5450 0.4300 0.7950 ;
      RECT 2.2950 1.6000 2.3850 1.9200 ;
      RECT 2.2950 1.5100 2.5500 1.6000 ;
      RECT 2.4600 0.7200 2.5500 1.5100 ;
      RECT 1.4500 0.6300 2.5500 0.7200 ;
      RECT 2.4300 0.4400 2.5500 0.6300 ;
      RECT 1.8950 0.4400 1.9850 0.6300 ;
      RECT 1.4500 0.7200 1.5450 1.0350 ;
  END
END OR6_X0P7M_A12TH

MACRO OR6_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.8600 0.3200 0.9500 0.6600 ;
        RECT 1.4150 0.3200 1.5050 0.6300 ;
        RECT 2.1250 0.3200 2.2150 0.5900 ;
        RECT 2.6450 0.3200 2.7350 0.5900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5500 1.0100 2.9450 1.1500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.7000 1.7550 1.9500 ;
        RECT 1.6500 0.6100 2.0050 0.7000 ;
        RECT 1.8350 0.4100 2.0050 0.6100 ;
    END
    ANTENNADIFFAREA 0.2534 ;
  END Y

  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0600 1.4500 1.3550 1.5500 ;
        RECT 1.2650 1.1050 1.3550 1.4500 ;
        RECT 1.1500 1.0050 1.3550 1.1050 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END F

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2150 1.2500 1.1550 1.3500 ;
        RECT 0.2150 1.1000 0.3050 1.2500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END E

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0400 0.9950 1.1500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END D

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2550 1.2400 3.1300 1.3500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0400 1.4500 3.3300 1.5500 ;
        RECT 3.2400 1.3200 3.3300 1.4500 ;
        RECT 2.0400 1.2950 2.1300 1.4500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.3950 1.8200 1.4850 2.0800 ;
        RECT 1.9250 1.8200 2.0150 2.0800 ;
        RECT 0.0800 1.7800 0.1700 2.0800 ;
        RECT 3.2300 1.7700 3.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6800 1.6400 1.5550 1.7300 ;
      RECT 1.4650 0.8800 1.5550 1.6400 ;
      RECT 0.6000 0.7900 1.5550 0.8800 ;
      RECT 0.6800 1.7300 0.8500 1.9300 ;
      RECT 0.6000 0.5400 0.6900 0.7900 ;
      RECT 1.1200 0.5400 1.2100 0.7900 ;
      RECT 2.5500 1.7300 2.7200 1.9500 ;
      RECT 1.8450 1.6400 2.7200 1.7300 ;
      RECT 1.8450 0.7900 2.9950 0.8800 ;
      RECT 2.9050 0.4700 2.9950 0.7900 ;
      RECT 1.8450 0.8800 1.9350 1.6400 ;
      RECT 2.3850 0.4700 2.4750 0.7900 ;
  END
END OR6_X1M_A12TH

MACRO OAI22_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7050 ;
        RECT 0.8750 0.3200 0.9650 0.7050 ;
        RECT 1.3950 0.3200 1.4850 0.7050 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3100 1.0500 0.8200 1.1600 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0800 1.0500 1.5500 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8450 1.0500 2.3550 1.1600 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5100 1.0500 2.9400 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.8950 3.1500 1.2500 ;
        RECT 0.0900 1.2500 3.3100 1.3500 ;
        RECT 1.8750 0.7950 3.1500 0.8950 ;
        RECT 0.0900 1.3500 0.1900 1.7000 ;
        RECT 0.6100 1.3500 0.7200 1.7000 ;
        RECT 2.6900 1.3500 2.7900 1.7200 ;
        RECT 3.2100 1.3500 3.3100 1.7200 ;
    END
    ANTENNADIFFAREA 1.0365 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 1.6550 1.7700 1.7450 2.0800 ;
        RECT 2.1750 1.7700 2.2650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6550 0.5900 3.3550 0.6800 ;
      RECT 0.0950 0.8000 1.7450 0.8900 ;
      RECT 1.6550 0.6800 1.7450 0.8000 ;
      RECT 0.0950 0.5000 0.1850 0.8000 ;
      RECT 0.8750 1.4600 1.4850 1.5500 ;
      RECT 1.3950 1.5500 1.4850 1.9250 ;
      RECT 0.3550 1.8250 0.9650 1.9150 ;
      RECT 0.8750 1.5500 0.9650 1.8250 ;
      RECT 0.3550 1.5150 0.4450 1.8250 ;
      RECT 2.4350 1.8300 3.0450 1.9200 ;
      RECT 2.9550 1.4900 3.0450 1.8300 ;
      RECT 1.9150 1.4550 2.5250 1.5450 ;
      RECT 2.4350 1.5450 2.5250 1.8300 ;
      RECT 1.9150 1.5450 2.0050 1.9350 ;
  END
END OAI22_X3M_A12TH

MACRO OAI22_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 2.5200 0.3200 2.6100 0.5800 ;
        RECT 3.0400 0.3200 3.1300 0.5800 ;
        RECT 3.5600 0.3200 3.6500 0.5800 ;
        RECT 4.0800 0.3200 4.1700 0.5800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 1.4500 3.9800 1.5500 ;
        RECT 0.6200 1.5500 0.7100 1.8800 ;
        RECT 1.6600 1.5500 1.7500 1.8800 ;
        RECT 2.8500 1.5500 2.9400 1.8800 ;
        RECT 3.8900 1.5500 3.9800 1.8800 ;
        RECT 2.2500 1.0200 2.3500 1.4500 ;
        RECT 2.0500 0.9300 2.3500 1.0200 ;
        RECT 2.0500 0.7500 2.1500 0.9300 ;
        RECT 0.4000 0.6600 2.1500 0.7500 ;
    END
    ANTENNADIFFAREA 1.2 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.0500 0.9050 1.1500 ;
        RECT 0.8150 0.9500 0.9050 1.0500 ;
        RECT 0.8150 0.8500 1.9150 0.9500 ;
        RECT 1.5450 0.9500 1.9150 0.9900 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6650 0.8500 4.0450 0.9500 ;
        RECT 2.6650 0.9500 3.0550 0.9950 ;
        RECT 3.6550 0.9500 4.0450 1.0050 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2950 1.2500 2.0550 1.3500 ;
        RECT 1.9650 1.2200 2.0550 1.2500 ;
        RECT 0.2950 1.1800 0.3850 1.2500 ;
        RECT 1.0250 1.1300 1.3950 1.2500 ;
        RECT 1.9650 1.1300 2.1550 1.2200 ;
        RECT 0.1750 1.0900 0.3850 1.1800 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4850 1.2500 4.3750 1.3500 ;
        RECT 3.2100 1.1100 3.5800 1.2500 ;
        RECT 2.4850 1.0900 2.5750 1.2500 ;
        RECT 4.2850 1.0900 4.3750 1.2500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1000 1.7700 0.1900 2.0800 ;
        RECT 1.1400 1.7700 1.2300 2.0800 ;
        RECT 2.3300 1.7700 2.4200 2.0800 ;
        RECT 3.3700 1.7700 3.4600 2.0800 ;
        RECT 4.4100 1.7700 4.5000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2600 0.6700 4.4700 0.7600 ;
      RECT 4.3000 0.4100 4.4700 0.6700 ;
      RECT 2.2600 0.7600 2.3500 0.7800 ;
      RECT 2.2600 0.5700 2.3500 0.6700 ;
      RECT 0.1800 0.4800 2.3500 0.5700 ;
      RECT 2.2600 0.4100 2.3500 0.4800 ;
      RECT 0.1800 0.5700 0.2700 0.8350 ;
      RECT 0.1800 0.4650 0.2700 0.4800 ;
      RECT 2.7400 0.4100 2.9100 0.6700 ;
      RECT 3.2600 0.4100 3.4300 0.6700 ;
      RECT 3.7800 0.4100 3.9500 0.6700 ;
  END
END OAI22_X4M_A12TH

MACRO OAI22_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 3.6400 0.3200 3.7300 0.4700 ;
        RECT 3.8900 0.3200 3.9800 0.4300 ;
        RECT 4.4100 0.3200 4.5000 0.5800 ;
        RECT 4.9300 0.3200 5.0200 0.5800 ;
        RECT 5.4500 0.3200 5.5400 0.5800 ;
        RECT 5.9700 0.3200 6.0600 0.5800 ;
    END
  END VSS

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1750 0.8500 3.0350 0.9500 ;
        RECT 0.1750 0.9500 0.2750 1.1900 ;
        RECT 0.8950 0.9500 1.2650 1.1500 ;
        RECT 1.9350 0.9500 2.3050 1.1500 ;
        RECT 2.9450 0.9500 3.0350 1.2300 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0050 0.9700 4.3750 1.1500 ;
        RECT 4.0050 0.9500 4.0950 0.9700 ;
        RECT 4.2850 0.9500 4.3750 0.9700 ;
        RECT 3.3050 0.8500 4.0950 0.9500 ;
        RECT 4.2850 0.8500 6.1350 0.9500 ;
        RECT 3.3050 0.9500 3.3950 1.2300 ;
        RECT 5.0450 0.9500 5.4150 1.1100 ;
        RECT 6.0450 0.9500 6.1350 1.1900 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3950 1.2500 2.4850 1.3500 ;
        RECT 2.3950 1.2000 2.4850 1.2500 ;
        RECT 0.3950 1.1100 0.7650 1.2500 ;
        RECT 1.4250 1.1100 1.7950 1.2500 ;
        RECT 2.3950 1.1100 2.8250 1.2000 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8250 1.2600 5.6550 1.3500 ;
        RECT 3.8250 1.2000 3.9150 1.2600 ;
        RECT 4.5250 1.2500 5.6550 1.2600 ;
        RECT 3.5050 1.1100 3.9150 1.2000 ;
        RECT 5.5650 1.2000 5.6550 1.2500 ;
        RECT 4.5250 1.1100 4.8950 1.2500 ;
        RECT 5.5650 1.1100 5.9350 1.2000 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5400 1.4500 5.8000 1.5500 ;
        RECT 0.5400 1.5500 0.6300 1.8800 ;
        RECT 1.5600 1.5500 1.6500 1.8800 ;
        RECT 2.6000 1.5500 2.6900 1.8800 ;
        RECT 3.6400 1.5500 3.7300 1.8800 ;
        RECT 4.6700 1.5500 4.7600 1.8800 ;
        RECT 5.7100 1.5500 5.8000 1.8800 ;
        RECT 3.1250 0.7500 3.2150 1.4500 ;
        RECT 0.7400 0.6600 3.2150 0.7500 ;
    END
    ANTENNADIFFAREA 1.802 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 1.0400 1.7700 1.1300 2.0800 ;
        RECT 2.0800 1.7700 2.1700 2.0800 ;
        RECT 3.1200 1.7700 3.2100 2.0800 ;
        RECT 4.1500 1.7700 4.2400 2.0800 ;
        RECT 5.1900 1.7700 5.2800 2.0800 ;
        RECT 6.2300 1.7700 6.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 6.2300 0.7600 6.3200 0.8200 ;
      RECT 3.3800 0.6700 6.3200 0.7600 ;
      RECT 6.2300 0.4100 6.3200 0.6700 ;
      RECT 3.3800 0.5700 3.4700 0.6650 ;
      RECT 0.4800 0.4800 3.4700 0.5700 ;
      RECT 3.3800 0.6650 4.2800 0.6700 ;
      RECT 4.1100 0.4100 4.2800 0.6650 ;
      RECT 4.6300 0.4100 4.8000 0.6700 ;
      RECT 5.1500 0.4100 5.3200 0.6700 ;
      RECT 5.6700 0.4100 5.8400 0.6700 ;
  END
END OAI22_X6M_A12TH

MACRO OAI22_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.6450 0.3200 ;
        RECT 4.7250 0.3200 4.8950 0.5800 ;
        RECT 5.0300 0.3200 5.1200 0.5800 ;
        RECT 5.5500 0.3200 5.6400 0.5800 ;
        RECT 6.0700 0.3200 6.1600 0.5800 ;
        RECT 6.5900 0.3200 6.6800 0.5800 ;
        RECT 7.1100 0.3200 7.2000 0.5800 ;
        RECT 7.6300 0.3200 7.7200 0.5800 ;
        RECT 8.1500 0.3200 8.2400 0.5800 ;
    END
  END VSS

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 0.8500 4.1600 0.9500 ;
        RECT 0.1900 0.9500 0.2800 1.1900 ;
        RECT 0.9800 0.9500 1.3500 1.0600 ;
        RECT 2.0200 0.9500 2.3900 1.0600 ;
        RECT 3.0400 0.9500 3.4100 1.0400 ;
        RECT 4.0700 0.9500 4.1600 1.1900 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.2500 3.9300 1.3500 ;
        RECT 3.5600 1.1200 3.9300 1.2500 ;
        RECT 0.4100 1.1100 0.8300 1.2500 ;
        RECT 1.5000 1.1100 1.8700 1.2500 ;
        RECT 2.5500 1.1100 2.9200 1.2500 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.2500 8.0950 1.3500 ;
        RECT 7.7250 1.1300 8.0950 1.2500 ;
        RECT 4.6500 1.1200 5.0200 1.2500 ;
        RECT 5.6450 1.1200 6.0150 1.2500 ;
        RECT 6.7350 1.1200 7.1050 1.2500 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6050 1.4500 7.9800 1.5500 ;
        RECT 0.6050 1.5500 0.6950 1.8800 ;
        RECT 1.6450 1.5500 1.7350 1.8800 ;
        RECT 2.6850 1.5500 2.7750 1.8800 ;
        RECT 3.7250 1.5500 3.8150 1.8800 ;
        RECT 4.7700 1.5500 4.8600 1.8800 ;
        RECT 5.8100 1.5500 5.9000 1.8800 ;
        RECT 6.8500 1.5500 6.9400 1.8800 ;
        RECT 7.8900 1.5500 7.9800 1.8800 ;
        RECT 4.2500 0.7600 4.3400 1.4500 ;
        RECT 0.8250 0.6700 4.3400 0.7600 ;
    END
    ANTENNADIFFAREA 2.401 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.6450 2.7200 ;
        RECT 0.0850 1.7700 0.1750 2.0800 ;
        RECT 1.1250 1.7700 1.2150 2.0800 ;
        RECT 2.1650 1.7700 2.2550 2.0800 ;
        RECT 3.2050 1.7700 3.2950 2.0800 ;
        RECT 4.2500 1.7700 4.3400 2.0800 ;
        RECT 5.2900 1.7700 5.3800 2.0800 ;
        RECT 6.3300 1.7700 6.4200 2.0800 ;
        RECT 7.3700 1.7700 7.4600 2.0800 ;
        RECT 8.4100 1.7700 8.5000 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4300 0.8500 8.3300 0.9500 ;
        RECT 4.4300 0.9500 4.5200 1.1950 ;
        RECT 5.1400 0.9500 5.5100 1.0400 ;
        RECT 6.1650 0.9500 6.5350 1.0400 ;
        RECT 7.2350 0.9500 7.6050 1.0400 ;
        RECT 8.2400 0.9500 8.3300 1.1900 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A1
  OBS
    LAYER M1 ;
      RECT 8.4100 0.7600 8.5000 0.8000 ;
      RECT 4.5050 0.6700 8.5000 0.7600 ;
      RECT 8.4100 0.4100 8.5000 0.6700 ;
      RECT 4.5050 0.5700 4.5950 0.6700 ;
      RECT 0.5650 0.4800 4.5950 0.5700 ;
      RECT 5.2500 0.4100 5.4200 0.6700 ;
      RECT 5.7700 0.4100 5.9400 0.6700 ;
      RECT 6.2900 0.4100 6.4600 0.6700 ;
      RECT 6.8100 0.4100 6.9800 0.6700 ;
      RECT 7.3300 0.4100 7.5000 0.6700 ;
      RECT 7.8500 0.4100 8.0200 0.6700 ;
  END
END OAI22_X8M_A12TH

MACRO OAI2XB1_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1000 0.3200 0.1900 0.8800 ;
        RECT 0.7100 0.3200 0.8000 0.4400 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9550 0.3750 1.3000 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8150 0.7550 0.9500 1.1650 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0100 1.1500 1.4400 ;
    END
    ANTENNAGATEAREA 0.0321 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6000 1.3500 1.6500 ;
        RECT 0.8550 1.6500 1.3500 1.7500 ;
        RECT 1.2300 0.4100 1.3500 0.6000 ;
        RECT 0.8550 1.7500 1.0250 1.9900 ;
    END
    ANTENNADIFFAREA 0.150825 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.2300 1.8400 1.3200 2.0800 ;
        RECT 0.3750 1.7800 0.4650 2.0800 ;
        RECT 0.1000 1.3750 0.1900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3000 1.4350 0.6300 1.5250 ;
      RECT 0.5400 0.8200 0.6300 1.4350 ;
      RECT 0.3000 0.7300 0.6300 0.8200 ;
      RECT 0.4500 0.5300 1.0600 0.6200 ;
      RECT 0.9700 0.4100 1.0600 0.5300 ;
      RECT 0.4500 0.4100 0.5400 0.5300 ;
  END
END OAI2XB1_X0P5M_A12TH

MACRO OAI2XB1_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1800 0.8900 ;
        RECT 0.8800 0.3200 0.9800 0.6750 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1800 1.3600 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.1200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8700 1.5500 1.4900 ;
        RECT 1.1500 1.4900 1.5500 1.5900 ;
        RECT 1.4050 0.5000 1.5500 0.8700 ;
        RECT 1.1500 1.5900 1.2500 1.7000 ;
    END
    ANTENNADIFFAREA 0.179075 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 0.9750 1.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0453 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.3750 1.8000 1.4750 2.0800 ;
        RECT 0.6200 1.7250 0.7100 2.0800 ;
        RECT 0.0900 1.4800 0.1800 2.0800 ;
        RECT 1.3750 1.7000 1.5500 1.8000 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4550 1.2400 0.7200 1.4100 ;
      RECT 0.3100 1.5400 0.5450 1.6300 ;
      RECT 0.4550 1.4100 0.5450 1.5400 ;
      RECT 0.4550 1.0900 0.5450 1.2400 ;
      RECT 0.3500 1.0000 0.5450 1.0900 ;
      RECT 0.3500 0.6800 0.4400 1.0000 ;
      RECT 0.6250 0.7950 1.2350 0.8850 ;
      RECT 1.1450 0.4750 1.2350 0.7950 ;
      RECT 0.6250 0.4750 0.7150 0.7950 ;
  END
END OAI2XB1_X0P7M_A12TH

MACRO OAI2XB1_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8600 ;
        RECT 0.8750 0.3200 0.9650 0.6500 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9800 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0273 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.2500 1.0800 1.3500 ;
        RECT 0.9800 1.0000 1.0800 1.2500 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8500 1.5500 1.5000 ;
        RECT 1.1350 1.5000 1.5500 1.6000 ;
        RECT 1.4050 0.4400 1.5500 0.8500 ;
        RECT 1.1350 1.6000 1.2350 1.9350 ;
    END
    ANTENNADIFFAREA 0.25835 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2200 1.0050 1.3500 1.3650 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.4100 1.7900 1.5000 2.0800 ;
        RECT 0.6150 1.7700 0.7050 2.0800 ;
        RECT 0.0800 1.5600 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.9850 0.8250 1.0750 ;
      RECT 0.2800 1.5750 0.5450 1.6650 ;
      RECT 0.4550 1.0750 0.5450 1.5750 ;
      RECT 0.3400 0.6500 0.4300 0.9850 ;
      RECT 0.6150 0.7700 1.2250 0.8600 ;
      RECT 1.1350 0.4400 1.2250 0.7700 ;
      RECT 0.6150 0.4400 0.7050 0.7700 ;
  END
END OAI2XB1_X1M_A12TH

MACRO OAI2XB1_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8600 ;
        RECT 0.8550 0.3200 0.9450 0.6500 ;
        RECT 1.3750 0.3200 1.4650 0.6500 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1700 1.2500 0.5900 1.3500 ;
    END
    ANTENNAGATEAREA 0.0375 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9500 1.0350 1.3400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8050 1.9500 1.5000 ;
        RECT 1.1100 1.5000 2.1200 1.6000 ;
        RECT 1.8500 0.7050 2.1200 0.8050 ;
        RECT 1.1100 1.6000 1.2100 1.9350 ;
    END
    ANTENNADIFFAREA 0.28 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9700 2.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.6300 1.7000 1.7300 2.0800 ;
        RECT 0.5950 1.6650 0.6850 2.0800 ;
        RECT 2.2300 1.5500 2.3200 2.0800 ;
        RECT 0.0800 1.5100 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.3050 1.6200 1.3950 ;
      RECT 1.5300 1.0350 1.6200 1.3050 ;
      RECT 0.3400 1.4550 0.7900 1.5450 ;
      RECT 0.7000 1.3950 0.7900 1.4550 ;
      RECT 0.7000 1.1000 0.7900 1.3050 ;
      RECT 0.3400 1.0100 0.7900 1.1000 ;
      RECT 0.3400 1.5450 0.4300 1.9200 ;
      RECT 0.3400 0.7150 0.4300 1.0100 ;
      RECT 1.6350 0.4800 2.3200 0.5700 ;
      RECT 2.2300 0.5700 2.3200 0.8800 ;
      RECT 0.5950 0.8000 1.7250 0.8900 ;
      RECT 1.6350 0.5700 1.7250 0.8000 ;
      RECT 0.5950 0.4500 0.6850 0.8000 ;
      RECT 1.1150 0.4500 1.2050 0.8000 ;
  END
END OAI2XB1_X1P4M_A12TH

MACRO OAI2XB1_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8500 ;
        RECT 0.8500 0.3200 0.9400 0.6450 ;
        RECT 1.3850 0.3200 1.4750 0.6450 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9000 2.1800 1.2250 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1250 1.5000 2.0600 1.6000 ;
        RECT 1.8500 0.7850 1.9500 1.5000 ;
        RECT 1.1250 1.6000 1.2150 1.9300 ;
        RECT 1.9600 1.6000 2.0600 1.7650 ;
        RECT 1.8500 0.6850 2.1100 0.7850 ;
    END
    ANTENNADIFFAREA 0.40865 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.5900 1.7700 0.6800 2.0800 ;
        RECT 1.6450 1.7700 1.7350 2.0800 ;
        RECT 0.0800 1.5100 0.1700 2.0800 ;
        RECT 2.2250 1.3400 2.3150 2.0800 ;
    END
  END VDD

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1150 1.2450 0.5350 1.3550 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9400 1.0500 1.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.6550 1.3000 1.6300 1.3900 ;
      RECT 1.5400 0.9650 1.6300 1.3000 ;
      RECT 0.3400 1.5050 0.7450 1.5950 ;
      RECT 0.6550 1.3900 0.7450 1.5050 ;
      RECT 0.6550 1.1000 0.7450 1.3000 ;
      RECT 0.3400 1.0100 0.7450 1.1000 ;
      RECT 0.3400 1.5950 0.4300 1.9150 ;
      RECT 0.3400 0.4650 0.4300 1.0100 ;
      RECT 1.6500 0.4800 2.3150 0.5700 ;
      RECT 2.2250 0.5700 2.3150 0.6900 ;
      RECT 0.5900 0.7650 1.7400 0.8550 ;
      RECT 1.6500 0.5700 1.7400 0.7650 ;
      RECT 0.5900 0.4400 0.6800 0.7650 ;
      RECT 1.1100 0.4450 1.2000 0.7650 ;
  END
END OAI2XB1_X2M_A12TH

MACRO OAI2XB1_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1100 0.3200 0.2000 0.8000 ;
        RECT 0.9350 0.3200 1.0250 0.7100 ;
        RECT 1.4550 0.3200 1.5450 0.7100 ;
        RECT 1.9750 0.3200 2.0650 0.7100 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0150 0.1700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6350 1.0500 2.1450 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8500 2.5500 1.2500 ;
        RECT 1.7100 1.2500 2.8700 1.3500 ;
        RECT 2.4500 0.7500 3.1250 0.8500 ;
        RECT 1.7100 1.3500 1.8100 1.7000 ;
        RECT 2.2400 1.3500 2.3400 1.7200 ;
        RECT 2.7700 1.3500 2.8700 1.7200 ;
        RECT 3.0250 0.4400 3.1250 0.7500 ;
    END
    ANTENNADIFFAREA 0.64155 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.6750 1.7700 0.7650 2.0800 ;
        RECT 1.1950 1.7700 1.2850 2.0800 ;
        RECT 0.1100 1.6100 0.2000 2.0800 ;
        RECT 2.5100 1.5550 2.6000 2.0800 ;
        RECT 3.0300 1.3550 3.1200 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6700 1.0500 3.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.1917 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 2.2350 0.4800 2.9200 0.5700 ;
      RECT 0.6750 0.8300 2.3250 0.9200 ;
      RECT 2.2350 0.5700 2.3250 0.8300 ;
      RECT 0.6750 0.4900 0.7650 0.8300 ;
      RECT 1.1950 0.4900 1.2850 0.8300 ;
      RECT 1.7150 0.4900 1.8050 0.8300 ;
      RECT 0.4550 1.0500 1.3650 1.1500 ;
      RECT 0.3700 1.3250 0.5450 1.7550 ;
      RECT 0.4550 1.1500 0.5450 1.3250 ;
      RECT 0.4550 0.9150 0.5450 1.0500 ;
      RECT 0.3700 0.4850 0.5450 0.9150 ;
      RECT 1.4550 1.8300 2.0650 1.9200 ;
      RECT 1.9750 1.5050 2.0650 1.8300 ;
      RECT 0.9350 1.5000 1.5450 1.5900 ;
      RECT 1.4550 1.5900 1.5450 1.8300 ;
      RECT 0.9350 1.5900 1.0250 1.9350 ;
  END
END OAI2XB1_X3M_A12TH

MACRO OAI2XB1_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.1100 0.3200 0.2000 0.6850 ;
        RECT 0.9550 0.3200 1.0450 0.7100 ;
        RECT 1.4750 0.3200 1.5650 0.7100 ;
        RECT 1.9950 0.3200 2.0850 0.7100 ;
        RECT 2.5150 0.3200 2.6050 0.7100 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1900 1.3100 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9300 1.0400 2.6600 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9950 1.2500 3.6500 1.3500 ;
        RECT 1.9950 1.3500 2.0850 1.7000 ;
        RECT 2.5150 1.3500 2.6050 1.7000 ;
        RECT 3.0300 1.3500 3.1300 1.7200 ;
        RECT 3.5500 1.3500 3.6500 1.7200 ;
        RECT 3.0300 0.7900 3.1300 1.2500 ;
        RECT 3.0300 0.6900 3.7150 0.7900 ;
    END
    ANTENNADIFFAREA 0.8286 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.1100 1.7700 0.2000 2.0800 ;
        RECT 0.9550 1.7700 1.0450 2.0800 ;
        RECT 1.4750 1.7700 1.5650 2.0800 ;
        RECT 3.2950 1.4950 3.3850 2.0800 ;
        RECT 3.8200 1.4950 3.9100 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.0500 3.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2559 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.3700 1.0500 1.4900 1.1500 ;
      RECT 0.3700 1.1500 0.4600 1.7200 ;
      RECT 0.3700 0.5400 0.4600 1.0500 ;
      RECT 1.7350 1.8300 2.8650 1.9200 ;
      RECT 2.7750 1.4900 2.8650 1.8300 ;
      RECT 0.6950 1.5000 1.8250 1.5900 ;
      RECT 1.7350 1.5900 1.8250 1.8300 ;
      RECT 2.2550 1.4900 2.3450 1.8300 ;
      RECT 0.6950 1.5900 0.7850 1.9300 ;
      RECT 1.2150 1.5900 1.3050 1.9300 ;
      RECT 2.7750 0.4800 3.9200 0.5700 ;
      RECT 3.8300 0.5700 3.9200 0.8900 ;
      RECT 0.6950 0.8300 2.8650 0.9200 ;
      RECT 2.7750 0.5700 2.8650 0.8300 ;
      RECT 0.6950 0.4600 0.7850 0.8300 ;
      RECT 1.2150 0.4600 1.3050 0.8300 ;
      RECT 1.7350 0.4600 1.8250 0.8300 ;
      RECT 2.2550 0.4600 2.3450 0.8300 ;
  END
END OAI2XB1_X4M_A12TH

MACRO OAI2XB1_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 1.8000 0.3200 1.9700 0.5750 ;
        RECT 2.0900 0.3200 2.1800 0.5800 ;
        RECT 2.6100 0.3200 2.7000 0.5800 ;
        RECT 3.1300 0.3200 3.2200 0.5800 ;
        RECT 3.6500 0.3200 3.7400 0.5800 ;
        RECT 4.1700 0.3200 4.2600 0.5800 ;
        RECT 4.6850 0.3200 4.7750 0.7350 ;
        RECT 5.2050 0.3200 5.2950 0.8050 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.0500 1.1000 1.1500 ;
    END
    ANTENNAGATEAREA 0.3846 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7150 1.0500 2.0850 1.1500 ;
        RECT 1.9950 0.9500 2.0850 1.0500 ;
        RECT 1.9950 0.8500 3.7950 0.9500 ;
        RECT 3.7050 0.9500 3.7950 1.0600 ;
        RECT 2.7350 0.9500 3.1050 1.1500 ;
        RECT 3.7050 1.0600 4.1350 1.1500 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A0

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8100 1.0500 5.2300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1482 ;
  END A1N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1300 1.4500 4.0000 1.5500 ;
        RECT 0.6100 1.5500 0.7000 1.8800 ;
        RECT 1.1300 1.5500 1.2200 1.8800 ;
        RECT 1.8600 1.5500 1.9500 1.8800 ;
        RECT 2.8700 1.5500 2.9600 1.8800 ;
        RECT 3.9100 1.5500 4.0000 1.8800 ;
        RECT 0.1300 0.9600 0.2200 1.4500 ;
        RECT 0.1300 0.8700 1.3000 0.9600 ;
        RECT 0.6100 0.6600 0.7800 0.8700 ;
        RECT 1.1300 0.6600 1.3000 0.8700 ;
        RECT 0.1300 0.5350 0.2200 0.8700 ;
    END
    ANTENNADIFFAREA 1.2438 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 1.4000 1.7700 1.4900 2.0800 ;
        RECT 2.3500 1.7700 2.4400 2.0800 ;
        RECT 3.3900 1.7700 3.4800 2.0800 ;
        RECT 4.3700 1.7700 4.4600 2.0800 ;
        RECT 0.3500 1.6550 0.4400 2.0800 ;
        RECT 0.8700 1.6550 0.9600 2.0800 ;
        RECT 4.6850 1.6200 4.7750 2.0800 ;
        RECT 5.2050 1.6200 5.2950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.4500 0.6700 4.5600 0.7600 ;
      RECT 4.4300 0.6650 4.5600 0.6700 ;
      RECT 4.4300 0.4250 4.5200 0.6650 ;
      RECT 1.4500 0.5700 1.5900 0.6700 ;
      RECT 0.3900 0.4800 1.5900 0.5700 ;
      RECT 1.5000 0.4250 1.5900 0.4800 ;
      RECT 0.3900 0.5700 0.4800 0.7800 ;
      RECT 0.3900 0.4100 0.4800 0.4800 ;
      RECT 0.9100 0.5700 1.0000 0.7800 ;
      RECT 0.9100 0.4100 1.0000 0.4800 ;
      RECT 2.3500 0.4250 2.4400 0.6700 ;
      RECT 2.8700 0.4250 2.9600 0.6700 ;
      RECT 3.3900 0.4250 3.4800 0.6700 ;
      RECT 3.9100 0.4250 4.0000 0.6700 ;
      RECT 1.5050 1.0000 1.5950 1.2400 ;
      RECT 1.5050 1.2400 5.0350 1.3300 ;
      RECT 4.2700 1.0100 4.3600 1.2400 ;
      RECT 4.6100 0.8700 5.0350 0.9600 ;
      RECT 4.6100 0.9600 4.7000 1.2400 ;
      RECT 4.9450 1.3300 5.0350 1.6350 ;
      RECT 4.9450 0.4900 5.0350 0.8700 ;
      RECT 2.2050 1.0700 2.5750 1.3300 ;
      RECT 3.2450 1.0700 3.6150 1.3300 ;
  END
END OAI2XB1_X6M_A12TH

MACRO OAI2XB1_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 2.1600 0.3200 2.2500 0.6350 ;
        RECT 2.6800 0.3200 2.7700 0.6350 ;
        RECT 3.2000 0.3200 3.2900 0.6350 ;
        RECT 3.7200 0.3200 3.8100 0.6350 ;
        RECT 4.2400 0.3200 4.3300 0.6350 ;
        RECT 4.7600 0.3200 4.8500 0.6350 ;
        RECT 5.2800 0.3200 5.3700 0.6350 ;
        RECT 5.8000 0.3200 5.8900 0.6350 ;
        RECT 6.3100 0.3200 6.4000 0.6350 ;
        RECT 6.8300 0.3200 6.9200 0.6350 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 1.2500 1.7350 1.3500 ;
    END
    ANTENNAGATEAREA 0.5124 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2850 1.0400 2.6800 1.1500 ;
        RECT 2.5900 0.9950 2.6800 1.0400 ;
        RECT 2.5900 0.9050 5.7350 0.9950 ;
        RECT 3.3150 0.9950 3.6850 1.1500 ;
        RECT 4.3650 0.9950 4.7350 1.1500 ;
        RECT 5.3650 0.9950 5.7350 1.1400 ;
    END
    ANTENNAGATEAREA 0.72 ;
  END A0

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4400 1.0500 6.8600 1.1500 ;
    END
    ANTENNAGATEAREA 0.195 ;
  END A1N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4500 5.6200 1.5500 ;
        RECT 0.1600 1.5500 0.2500 1.8800 ;
        RECT 0.6800 1.5500 0.7700 1.8800 ;
        RECT 1.2000 1.5500 1.2900 1.8800 ;
        RECT 1.7200 1.5500 1.8100 1.8800 ;
        RECT 2.4400 1.5500 2.5300 1.8800 ;
        RECT 3.4600 1.5500 3.5500 1.8800 ;
        RECT 4.5000 1.5500 4.5900 1.8800 ;
        RECT 5.5300 1.5500 5.6200 1.8800 ;
        RECT 0.0800 1.0400 0.1700 1.4500 ;
        RECT 0.0800 0.9500 1.6900 1.0400 ;
        RECT 0.5600 0.6600 0.7300 0.9500 ;
        RECT 1.0800 0.6600 1.2500 0.9500 ;
        RECT 1.6000 0.6600 1.7700 0.9500 ;
        RECT 0.0800 0.6050 0.1700 0.9500 ;
    END
    ANTENNADIFFAREA 1.6643 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 2.9400 1.7700 3.0300 2.0800 ;
        RECT 3.9800 1.7700 4.0700 2.0800 ;
        RECT 5.0200 1.7700 5.1100 2.0800 ;
        RECT 6.0000 1.7700 6.0900 2.0800 ;
        RECT 6.3100 1.7700 6.4000 2.0800 ;
        RECT 6.8300 1.7700 6.9200 2.0800 ;
        RECT 0.4200 1.6400 0.5100 2.0800 ;
        RECT 0.9400 1.6400 1.0300 2.0800 ;
        RECT 1.4600 1.6400 1.5500 2.0800 ;
        RECT 1.9800 1.6400 2.0700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.9000 0.7250 6.1500 0.8150 ;
      RECT 6.0600 0.4450 6.1500 0.7250 ;
      RECT 1.9000 0.8150 1.9900 0.8300 ;
      RECT 1.9000 0.5700 1.9900 0.7250 ;
      RECT 0.3400 0.4800 1.9900 0.5700 ;
      RECT 1.9000 0.4600 1.9900 0.4800 ;
      RECT 0.3400 0.5700 0.4300 0.8500 ;
      RECT 0.8600 0.5700 0.9500 0.8500 ;
      RECT 1.3800 0.5700 1.4700 0.8500 ;
      RECT 2.4200 0.4450 2.5100 0.7250 ;
      RECT 2.9400 0.4450 3.0300 0.7250 ;
      RECT 3.4600 0.4450 3.5500 0.7250 ;
      RECT 3.9800 0.4450 4.0700 0.7250 ;
      RECT 4.5000 0.4450 4.5900 0.7250 ;
      RECT 5.0200 0.4450 5.1100 0.7250 ;
      RECT 5.5400 0.4450 5.6300 0.7250 ;
      RECT 2.0850 1.2500 6.6600 1.3500 ;
      RECT 2.0850 1.0000 2.1750 1.2500 ;
      RECT 5.9050 1.0000 5.9950 1.2500 ;
      RECT 6.2400 0.9600 6.3300 1.2500 ;
      RECT 6.2400 0.8700 6.6600 0.9600 ;
      RECT 6.5700 1.3500 6.6600 1.7200 ;
      RECT 6.5700 0.4900 6.6600 0.8700 ;
      RECT 2.7950 1.0850 3.1650 1.3500 ;
      RECT 3.8350 1.0850 4.2050 1.3500 ;
      RECT 4.8550 1.1300 5.2250 1.3500 ;
  END
END OAI2XB1_X8M_A12TH

MACRO OAI31_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.5500 ;
        RECT 0.5850 0.3200 0.7750 0.4650 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7350 0.5600 1.1900 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9950 0.7450 1.1500 1.1600 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END B0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 0.7450 0.3600 1.1600 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7450 0.8350 1.1600 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8550 1.4550 1.3500 1.5550 ;
        RECT 0.8550 1.5550 1.0250 1.9050 ;
        RECT 1.2500 0.5300 1.3500 1.4550 ;
        RECT 1.1000 0.4300 1.3500 0.5300 ;
    END
    ANTENNADIFFAREA 0.1111 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0550 1.8450 0.2250 2.0800 ;
        RECT 1.1150 1.7750 1.2850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3500 0.5550 0.9900 0.6450 ;
      RECT 0.8900 0.4100 0.9900 0.5550 ;
      RECT 0.3500 0.4100 0.4500 0.5550 ;
  END
END OAI31_X0P5M_A12TH

MACRO OAI31_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.5000 ;
        RECT 0.5850 0.3200 0.7750 0.3850 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7000 0.5600 1.1900 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9950 0.7450 1.1500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0297 ;
  END B0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 0.7450 0.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7450 0.8350 1.1500 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8550 1.4450 1.3500 1.5450 ;
        RECT 0.8550 1.5450 1.0250 1.7500 ;
        RECT 1.2500 0.5450 1.3500 1.4450 ;
        RECT 1.1000 0.4450 1.3500 0.5450 ;
    END
    ANTENNADIFFAREA 0.15725 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0550 1.8450 0.2250 2.0800 ;
        RECT 1.1150 1.6700 1.2850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3500 0.4900 0.9900 0.5800 ;
      RECT 0.3500 0.4100 0.4500 0.4900 ;
      RECT 0.8900 0.4100 0.9900 0.4900 ;
  END
END OAI31_X0P7M_A12TH

MACRO OAI31_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.4450 ;
        RECT 0.5850 0.3200 0.7750 0.3800 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7000 0.5500 1.1900 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9950 0.7450 1.1500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0423 ;
  END B0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 0.7450 0.3600 1.1900 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7450 0.8350 1.1150 ;
        RECT 0.6500 1.1150 0.7500 1.2200 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8550 1.6500 1.3500 1.7500 ;
        RECT 0.8550 1.7500 1.0250 1.9900 ;
        RECT 1.2500 0.5500 1.3500 1.6500 ;
        RECT 1.1000 0.4500 1.3500 0.5500 ;
    END
    ANTENNADIFFAREA 0.22245 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1500 1.9450 1.2500 2.0800 ;
        RECT 0.0550 1.8450 0.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3500 0.4900 0.9900 0.5800 ;
      RECT 0.3500 0.4100 0.4500 0.4900 ;
      RECT 0.8900 0.4100 0.9900 0.4900 ;
  END
END OAI31_X1M_A12TH

MACRO OAI31_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.6050 2.0300 1.7800 2.0800 ;
        RECT 0.0450 1.8450 0.2250 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.8600 0.3200 0.9600 0.7600 ;
        RECT 1.3450 0.3200 1.5150 0.5100 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0400 0.9800 2.1550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0597 ;
  END B0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1300 0.8500 1.6350 0.9500 ;
        RECT 1.5300 0.9500 1.6350 1.2050 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.1000 1.1550 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.4500 1.3750 1.5500 ;
        RECT 0.4500 1.2450 0.5500 1.4500 ;
        RECT 1.2500 1.0500 1.3750 1.4500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8250 1.9500 1.6500 ;
        RECT 0.8250 1.6500 2.0000 1.7500 ;
        RECT 1.8500 0.7250 2.0000 0.8250 ;
        RECT 0.8250 1.7500 0.9950 1.9500 ;
        RECT 1.9000 1.7500 2.0000 1.9650 ;
        RECT 1.9000 0.4250 2.0000 0.7250 ;
    END
    ANTENNADIFFAREA 0.30535 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.0700 0.6100 1.7350 0.7000 ;
      RECT 1.6450 0.4800 1.7350 0.6100 ;
  END
END OAI31_X1P4M_A12TH

MACRO OAI31_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3000 0.3200 0.4850 0.5100 ;
        RECT 0.8150 0.3200 1.0050 0.5100 ;
        RECT 1.3450 0.3200 1.5150 0.5100 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9800 2.1550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END B0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1850 0.8500 1.6350 0.9400 ;
        RECT 0.1850 0.9400 0.3500 1.1900 ;
        RECT 1.5300 0.9400 1.6350 1.1000 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.1000 1.1550 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.4500 1.3750 1.5500 ;
        RECT 0.4500 1.0500 0.5500 1.4500 ;
        RECT 1.2500 1.0500 1.3750 1.4500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.7700 1.9500 1.6500 ;
        RECT 0.8250 1.6500 2.0350 1.7500 ;
        RECT 1.8500 0.6700 2.0350 0.7700 ;
        RECT 0.8250 1.7500 0.9950 1.9500 ;
        RECT 1.8650 1.7500 2.0350 1.9900 ;
    END
    ANTENNADIFFAREA 0.323 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.6050 2.0300 1.7800 2.0800 ;
        RECT 2.1600 2.0000 2.2600 2.0800 ;
        RECT 0.0450 1.8450 0.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6050 0.4800 2.2950 0.5800 ;
      RECT 0.0800 0.6100 1.6950 0.7000 ;
      RECT 1.6050 0.5800 1.6950 0.6100 ;
      RECT 0.0800 0.5100 0.1800 0.6100 ;
  END
END OAI31_X2M_A12TH

MACRO OAI31_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.5400 ;
        RECT 0.8350 0.3200 1.0050 0.5400 ;
        RECT 1.3550 0.3200 1.5250 0.5350 ;
        RECT 1.8750 0.3200 2.0450 0.5350 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8500 2.3500 0.9500 ;
        RECT 1.6500 0.9500 1.7500 1.0500 ;
        RECT 2.2500 0.9500 2.3500 1.1600 ;
        RECT 1.3300 1.0500 1.7500 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.5500 2.5500 1.9400 ;
        RECT 2.4500 1.5400 3.1450 1.5500 ;
        RECT 2.9700 1.5500 3.0700 1.9400 ;
        RECT 1.3550 1.4400 3.1450 1.5400 ;
        RECT 1.3550 1.5400 1.5250 1.7300 ;
        RECT 3.0450 0.7600 3.1450 1.4400 ;
        RECT 2.5550 0.6600 3.1450 0.7600 ;
    END
    ANTENNADIFFAREA 0.553 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4800 1.0500 2.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.1266 ;
  END B0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 0.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.2500 1.9500 1.3500 ;
        RECT 1.8500 1.1500 1.9500 1.2500 ;
        RECT 1.0500 1.0400 1.1500 1.2500 ;
        RECT 1.8500 1.0500 2.0800 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0550 1.8450 0.2250 2.0800 ;
        RECT 0.5750 1.8450 0.7450 2.0800 ;
        RECT 2.6750 1.8400 2.8450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8350 1.8300 2.0450 1.9200 ;
      RECT 1.8750 1.6300 2.0450 1.8300 ;
      RECT 0.8350 1.9200 1.0050 1.9650 ;
      RECT 0.8350 1.7550 1.0050 1.8300 ;
      RECT 0.3150 1.6650 1.0050 1.7550 ;
      RECT 0.3150 1.7550 0.4850 1.9650 ;
      RECT 2.1900 0.4800 3.0250 0.5700 ;
      RECT 0.5750 0.6500 2.3600 0.7400 ;
      RECT 2.1900 0.5700 2.3600 0.6500 ;
      RECT 2.1900 0.4300 2.3600 0.4800 ;
      RECT 0.5750 0.4300 0.7450 0.6500 ;
      RECT 1.0950 0.4300 1.2650 0.6500 ;
      RECT 1.6150 0.4300 1.7850 0.6500 ;
  END
END OAI31_X3M_A12TH

MACRO OAI31_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.5900 0.3200 0.7600 0.4800 ;
        RECT 1.1100 0.3200 1.2800 0.4800 ;
        RECT 1.6300 0.3200 1.8000 0.4750 ;
        RECT 2.1500 0.3200 2.3200 0.4750 ;
        RECT 2.6800 0.3200 2.8500 0.4750 ;
        RECT 3.0050 0.3200 3.1750 0.4750 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 1.0350 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5550 1.0500 4.1200 1.1500 ;
    END
    ANTENNAGATEAREA 0.1683 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6300 1.4400 4.3500 1.5400 ;
        RECT 3.7050 1.5400 4.3500 1.5500 ;
        RECT 1.6300 1.5400 1.8000 1.7300 ;
        RECT 2.6700 1.5400 2.8400 1.7300 ;
        RECT 4.2500 0.7600 4.3500 1.4400 ;
        RECT 4.2500 1.5500 4.3500 1.7650 ;
        RECT 3.7050 1.5500 3.8050 1.9750 ;
        RECT 3.5450 0.6600 4.3500 0.7600 ;
        RECT 4.2250 1.7650 4.3500 1.9750 ;
        RECT 4.1050 0.4250 4.2050 0.6600 ;
    END
    ANTENNADIFFAREA 0.724 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9250 0.8500 2.6250 0.9500 ;
        RECT 1.9250 0.9500 2.0250 1.0500 ;
        RECT 2.5250 0.9500 2.6250 1.0450 ;
        RECT 1.6050 1.0500 2.0250 1.1500 ;
        RECT 2.5250 1.0450 2.8500 1.1450 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2250 1.2600 3.2200 1.3500 ;
        RECT 1.2250 1.2500 2.2250 1.2600 ;
        RECT 3.1200 1.0000 3.2200 1.2600 ;
        RECT 2.1250 1.1500 2.2250 1.2500 ;
        RECT 1.2250 1.0400 1.3500 1.2500 ;
        RECT 2.1250 1.0500 2.3550 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 3.4050 2.0400 3.5850 2.0800 ;
        RECT 0.3300 1.8450 0.5000 2.0800 ;
        RECT 0.8500 1.8450 1.0200 2.0800 ;
        RECT 3.9300 1.8450 4.1000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1100 1.8300 3.3450 1.9200 ;
      RECT 3.1600 1.6300 3.3450 1.8300 ;
      RECT 1.1100 1.9200 1.2800 1.9650 ;
      RECT 1.1100 1.7550 1.2800 1.8300 ;
      RECT 0.0700 1.6650 1.2800 1.7550 ;
      RECT 2.1500 1.6300 2.3200 1.8300 ;
      RECT 0.0700 1.7550 0.2400 1.9650 ;
      RECT 0.5900 1.7550 0.7600 1.9650 ;
      RECT 3.2650 0.4800 3.9950 0.5700 ;
      RECT 0.3250 0.6500 3.4350 0.7400 ;
      RECT 3.2650 0.5700 3.4350 0.6500 ;
      RECT 3.2650 0.4300 3.4350 0.4800 ;
      RECT 0.3250 0.4300 0.5000 0.6500 ;
      RECT 0.8500 0.4300 1.0200 0.6500 ;
      RECT 1.3700 0.4300 1.5400 0.6500 ;
      RECT 1.8900 0.4300 2.0600 0.6500 ;
      RECT 2.4100 0.4300 2.5800 0.6500 ;
  END
END OAI31_X4M_A12TH

MACRO OAI31_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.5650 0.3200 0.7350 0.4800 ;
        RECT 1.0850 0.3200 1.2550 0.4800 ;
        RECT 1.6050 0.3200 1.7750 0.4800 ;
        RECT 2.1250 0.3200 2.2950 0.4750 ;
        RECT 2.6450 0.3200 2.8150 0.4750 ;
        RECT 3.1650 0.3200 3.3350 0.4750 ;
        RECT 3.6850 0.3200 3.8550 0.4750 ;
        RECT 4.2050 0.3200 4.3750 0.4750 ;
        RECT 4.5900 0.3200 4.7600 0.4750 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 1.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.4686 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1000 1.0500 6.1000 1.1500 ;
    END
    ANTENNAGATEAREA 0.2535 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1250 1.4400 6.4550 1.5400 ;
        RECT 5.2900 1.5400 6.4550 1.5500 ;
        RECT 2.1250 1.5400 2.2950 1.7300 ;
        RECT 3.1650 1.5400 3.3350 1.7300 ;
        RECT 4.2050 1.5400 4.3750 1.7300 ;
        RECT 6.3550 0.7600 6.4550 1.4400 ;
        RECT 5.2900 1.5500 5.3900 1.9900 ;
        RECT 5.8100 1.5500 5.9100 1.9900 ;
        RECT 6.3300 1.5500 6.4550 1.9900 ;
        RECT 5.1300 0.6600 6.4550 0.7600 ;
        RECT 6.2100 0.4250 6.3100 0.6600 ;
    END
    ANTENNADIFFAREA 1.040325 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.8500 4.1450 0.9500 ;
        RECT 2.2500 0.9500 2.3500 1.0500 ;
        RECT 3.0500 0.9500 3.1500 1.0500 ;
        RECT 4.0450 0.9500 4.1450 1.0500 ;
        RECT 2.1000 1.0500 2.3500 1.1500 ;
        RECT 3.0500 1.0500 3.3500 1.1500 ;
        RECT 4.0450 1.0500 4.3950 1.1500 ;
    END
    ANTENNAGATEAREA 0.4686 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 4.9900 2.0400 5.1700 2.0800 ;
        RECT 0.3050 1.8450 0.4750 2.0800 ;
        RECT 0.8250 1.8450 0.9950 2.0800 ;
        RECT 1.3450 1.8450 1.5150 2.0800 ;
        RECT 5.5150 1.8450 5.6850 2.0800 ;
        RECT 6.0350 1.8450 6.2050 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7200 1.2500 4.8050 1.3500 ;
        RECT 2.6200 1.1500 2.7200 1.2500 ;
        RECT 3.6500 1.1500 3.7500 1.2500 ;
        RECT 1.7200 1.0400 1.8450 1.2500 ;
        RECT 4.7050 1.0000 4.8050 1.2500 ;
        RECT 2.6200 1.0500 2.8500 1.1500 ;
        RECT 3.6500 1.0500 3.8700 1.1500 ;
    END
    ANTENNAGATEAREA 0.4686 ;
  END A1
  OBS
    LAYER M1 ;
      RECT 1.6050 1.8300 4.9300 1.9200 ;
      RECT 4.7450 1.6300 4.9300 1.8300 ;
      RECT 1.6050 1.9200 1.7750 1.9650 ;
      RECT 1.6050 1.7550 1.7750 1.8300 ;
      RECT 0.0450 1.6650 1.7750 1.7550 ;
      RECT 2.6450 1.6300 2.8150 1.8300 ;
      RECT 3.6850 1.6300 3.8550 1.8300 ;
      RECT 0.0450 1.7550 0.2150 1.9650 ;
      RECT 0.5650 1.7550 0.7350 1.9650 ;
      RECT 1.0850 1.7550 1.2550 1.9650 ;
      RECT 4.8500 0.4800 6.0950 0.5700 ;
      RECT 0.3050 0.6500 5.0200 0.7400 ;
      RECT 4.8500 0.5700 5.0200 0.6500 ;
      RECT 4.8500 0.4300 5.0200 0.4800 ;
      RECT 0.3050 0.4300 0.4750 0.6500 ;
      RECT 0.8250 0.4300 0.9950 0.6500 ;
      RECT 1.3450 0.4300 1.5150 0.6500 ;
      RECT 1.8650 0.4300 2.0350 0.6500 ;
      RECT 2.3850 0.4300 2.5550 0.6500 ;
      RECT 2.9050 0.4300 3.0750 0.6500 ;
      RECT 3.4250 0.4300 3.5950 0.6500 ;
      RECT 3.9450 0.4300 4.1150 0.6500 ;
  END
END OAI31_X6M_A12TH

MACRO OR2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7400 ;
        RECT 0.6700 0.3200 0.7700 0.7150 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.6350 1.7400 0.8050 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7150 1.1500 1.6000 ;
        RECT 0.9500 1.6000 1.1500 1.7000 ;
        RECT 0.8950 0.6150 1.1500 0.7150 ;
        RECT 0.9500 1.7000 1.0500 1.9800 ;
        RECT 0.8950 0.4100 1.0650 0.6150 ;
    END
    ANTENNADIFFAREA 0.17845 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0100 0.5500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9950 0.1600 1.4150 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0900 1.5250 0.8400 1.6150 ;
      RECT 0.7500 0.9000 0.8400 1.5250 ;
      RECT 0.3550 0.8100 0.8400 0.9000 ;
      RECT 0.3550 0.5300 0.4450 0.8100 ;
      RECT 0.0900 1.6150 0.1800 1.9800 ;
  END
END OR2_X0P5M_A12TH

MACRO OR2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7450 ;
        RECT 0.6900 0.3200 0.7900 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.6150 1.7350 0.7850 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7300 1.1500 1.4500 ;
        RECT 0.9750 1.4500 1.1500 1.5500 ;
        RECT 0.9150 0.6300 1.1500 0.7300 ;
        RECT 0.9750 1.5500 1.0750 1.8800 ;
        RECT 0.9150 0.4200 1.0850 0.6300 ;
    END
    ANTENNADIFFAREA 0.2529 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0100 0.5500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0399 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9950 0.1600 1.4150 ;
    END
    ANTENNAGATEAREA 0.0399 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0900 1.5250 0.8600 1.6150 ;
      RECT 0.7700 0.9000 0.8600 1.5250 ;
      RECT 0.3550 0.8100 0.8600 0.9000 ;
      RECT 0.3550 0.5300 0.4450 0.8100 ;
      RECT 0.0900 1.6150 0.1800 1.9800 ;
  END
END OR2_X0P7M_A12TH

MACRO OR2_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 1.8150 0.3200 1.9050 0.5800 ;
        RECT 2.3350 0.3200 2.4250 0.5800 ;
        RECT 2.8550 0.3200 2.9450 0.5800 ;
        RECT 3.3750 0.3200 3.4650 0.5800 ;
        RECT 3.9700 0.3200 4.0600 0.5800 ;
        RECT 4.4900 0.3200 4.5800 0.6500 ;
        RECT 5.0100 0.3200 5.1000 0.6500 ;
        RECT 5.5300 0.3200 5.6200 0.6500 ;
        RECT 6.0500 0.3200 6.1400 0.6500 ;
        RECT 6.5700 0.3200 6.6600 0.6500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7850 0.8500 3.8800 0.9500 ;
        RECT 0.7850 0.9500 1.2000 1.0400 ;
        RECT 1.8350 0.9500 2.0450 1.1500 ;
        RECT 2.7500 0.9500 3.1200 1.0650 ;
        RECT 3.7800 0.9500 3.8800 1.1700 ;
    END
    ANTENNAGATEAREA 0.5544 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.2500 3.6400 1.3500 ;
        RECT 0.4050 1.1800 0.7600 1.2500 ;
        RECT 2.2300 1.2300 3.6400 1.2500 ;
        RECT 1.3200 1.1600 1.6600 1.2500 ;
        RECT 2.2300 1.1200 2.6000 1.2300 ;
        RECT 3.2650 1.1200 3.6400 1.2300 ;
    END
    ANTENNAGATEAREA 0.5544 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2200 1.4200 6.9250 1.5800 ;
        RECT 4.2200 1.5800 4.3250 1.8500 ;
        RECT 4.7450 1.5800 4.8450 1.8250 ;
        RECT 5.2650 1.5800 5.3650 1.8250 ;
        RECT 5.7850 1.5800 5.8850 1.8250 ;
        RECT 6.3050 1.5800 6.4050 1.8250 ;
        RECT 6.8250 1.5800 6.9250 1.8500 ;
        RECT 6.6200 0.9800 6.7800 1.4200 ;
        RECT 4.2250 0.8200 6.9250 0.9800 ;
        RECT 4.2250 0.5050 4.3250 0.8200 ;
        RECT 4.7450 0.5050 4.8450 0.8200 ;
        RECT 5.2650 0.5050 5.3650 0.8200 ;
        RECT 5.7850 0.5050 5.8850 0.8200 ;
        RECT 6.3050 0.5050 6.4050 0.8200 ;
        RECT 6.8250 0.5050 6.9250 0.8200 ;
    END
    ANTENNADIFFAREA 1.885 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 4.4900 1.7700 4.5800 2.0800 ;
        RECT 5.0100 1.7700 5.1000 2.0800 ;
        RECT 5.5300 1.7700 5.6200 2.0800 ;
        RECT 6.0500 1.7700 6.1400 2.0800 ;
        RECT 6.5700 1.7700 6.6600 2.0800 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 0.9950 1.7500 1.0850 2.0800 ;
        RECT 1.8950 1.7500 1.9850 2.0800 ;
        RECT 2.9150 1.7500 3.0050 2.0800 ;
        RECT 3.9700 1.7500 4.0600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.9700 1.0700 6.4300 1.1600 ;
      RECT 0.5450 1.5900 0.6350 1.9350 ;
      RECT 1.4450 1.5900 1.5350 1.9350 ;
      RECT 2.0350 0.4600 2.2050 0.6700 ;
      RECT 2.3950 1.5900 2.4850 1.9350 ;
      RECT 2.5950 0.4300 2.6850 0.6700 ;
      RECT 3.1150 0.4300 3.2050 0.6700 ;
      RECT 3.4350 1.5900 3.5250 1.9300 ;
      RECT 3.6350 0.4300 3.7250 0.6700 ;
      RECT 0.5450 1.5000 4.0600 1.5900 ;
      RECT 3.9700 1.1600 4.0600 1.5000 ;
      RECT 3.9700 0.7600 4.0600 1.0700 ;
      RECT 2.0350 0.6700 4.0600 0.7600 ;
  END
END OR2_X11M_A12TH

MACRO OR2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.8750 ;
        RECT 0.6700 0.3200 0.7700 0.6200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.6400 1.7800 0.7400 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.4500 ;
        RECT 0.9350 1.4500 1.1500 1.5500 ;
        RECT 0.9300 0.8500 1.1500 0.9500 ;
        RECT 0.9350 1.5500 1.0350 1.9100 ;
        RECT 0.9300 0.4950 1.0300 0.8500 ;
    END
    ANTENNADIFFAREA 0.337675 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4400 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9950 0.1600 1.4150 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0850 1.5600 0.8100 1.6600 ;
      RECT 0.7100 0.8900 0.8100 1.5600 ;
      RECT 0.3500 0.7900 0.8100 0.8900 ;
      RECT 0.3500 0.6800 0.4500 0.7900 ;
      RECT 0.0850 1.6600 0.1850 1.9800 ;
  END
END OR2_X1M_A12TH

MACRO OR2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.6150 ;
        RECT 0.6850 0.3200 0.7850 0.7100 ;
        RECT 1.2050 0.3200 1.3050 0.7100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6400 1.7700 0.7400 2.0800 ;
        RECT 1.2050 1.7700 1.3050 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.4500 ;
        RECT 0.9450 1.4500 1.3500 1.5500 ;
        RECT 0.9450 0.8500 1.3500 0.9500 ;
        RECT 0.9450 1.5500 1.0450 1.9700 ;
        RECT 0.9450 0.4100 1.0450 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0100 0.5500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0714 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7600 0.1600 1.2000 ;
    END
    ANTENNAGATEAREA 0.0714 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0750 1.1250 1.1850 ;
      RECT 0.0950 1.5400 0.7900 1.6300 ;
      RECT 0.7000 1.1850 0.7900 1.5400 ;
      RECT 0.7000 0.9000 0.7900 1.0750 ;
      RECT 0.3550 0.8100 0.7900 0.9000 ;
      RECT 0.3550 0.4200 0.4450 0.8100 ;
      RECT 0.0950 1.6300 0.1850 1.9800 ;
  END
END OR2_X1P4M_A12TH

MACRO OAI21_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.5800 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9250 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9250 0.5600 1.3100 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8450 0.8050 0.9550 1.1900 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.6100 1.1500 1.3000 ;
        RECT 0.6500 1.3000 1.1500 1.4000 ;
        RECT 0.8900 0.5200 1.1500 0.6100 ;
        RECT 0.6500 1.4000 0.7500 1.7600 ;
    END
    ANTENNADIFFAREA 0.2731 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.1350 1.7700 0.2250 2.0800 ;
        RECT 0.9300 1.5550 1.0200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1350 0.7000 0.7450 0.8000 ;
      RECT 0.6550 0.4100 0.7450 0.7000 ;
      RECT 0.1350 0.4100 0.2250 0.7000 ;
  END
END OAI21_X1M_A12TH

MACRO OAI21_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3950 0.3200 0.4850 0.6600 ;
        RECT 0.9150 0.3200 1.0050 0.6600 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 1.1150 1.3500 ;
        RECT 1.0150 1.0200 1.1150 1.2500 ;
        RECT 0.2400 1.0000 0.3400 1.2500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4700 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2950 1.0500 1.7300 1.1500 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.7900 1.9500 1.2500 ;
        RECT 1.5050 1.2500 1.9500 1.3500 ;
        RECT 1.4400 0.6900 1.9500 0.7900 ;
        RECT 1.5050 1.3500 1.6050 1.4500 ;
        RECT 0.6550 1.4500 1.6050 1.5500 ;
        RECT 0.6550 1.5500 0.7450 1.8800 ;
    END
    ANTENNADIFFAREA 0.28 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.1750 1.7300 1.2650 2.0800 ;
        RECT 0.1350 1.5100 0.2250 2.0800 ;
        RECT 1.7700 1.4400 1.8600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.2150 0.4800 1.9150 0.5700 ;
      RECT 0.1350 0.7800 1.3050 0.8700 ;
      RECT 1.2150 0.5700 1.3050 0.7800 ;
      RECT 0.1350 0.6600 0.2250 0.7800 ;
      RECT 0.6550 0.6600 0.7450 0.7800 ;
  END
END OAI21_X1P4M_A12TH

MACRO OAI21_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3950 0.3200 0.4850 0.6700 ;
        RECT 0.9300 0.3200 1.0200 0.6700 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3600 1.0400 1.7500 1.1600 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 1.2000 1.3500 ;
        RECT 0.2400 0.9700 0.3550 1.2500 ;
        RECT 1.1000 0.9700 1.2000 1.2500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.7950 1.9500 1.3350 ;
        RECT 1.5200 1.3350 1.9500 1.4350 ;
        RECT 1.4600 0.6950 1.9500 0.7950 ;
        RECT 1.5200 1.4350 1.6200 1.4500 ;
        RECT 0.6700 1.4500 1.6200 1.5500 ;
        RECT 0.6700 1.5500 0.7600 1.8800 ;
        RECT 1.5200 1.5500 1.6200 1.7650 ;
    END
    ANTENNADIFFAREA 0.40865 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1350 1.7700 0.2250 2.0800 ;
        RECT 1.1900 1.7700 1.2800 2.0800 ;
        RECT 1.7850 1.5550 1.8750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1950 0.4800 1.9350 0.5700 ;
      RECT 0.1350 0.7600 1.2850 0.8500 ;
      RECT 1.1950 0.5700 1.2850 0.7600 ;
      RECT 0.1350 0.4200 0.2250 0.7600 ;
      RECT 0.6700 0.4200 0.7600 0.7600 ;
  END
END OAI21_X2M_A12TH

MACRO OAI21_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6450 ;
        RECT 0.8750 0.3200 0.9650 0.6450 ;
        RECT 1.3950 0.3200 1.4850 0.6450 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0700 1.0500 1.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0500 0.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8600 1.0500 2.3400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1917 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1300 1.2500 2.5500 1.3500 ;
        RECT 1.1300 1.3500 1.2300 1.7200 ;
        RECT 1.6600 1.3500 1.7500 1.7200 ;
        RECT 2.2500 1.3500 2.3400 1.7200 ;
        RECT 2.4500 0.9500 2.5500 1.2500 ;
        RECT 1.9500 0.8500 2.6000 0.9500 ;
        RECT 1.9500 0.6600 2.1200 0.8500 ;
        RECT 2.5100 0.4350 2.6000 0.8500 ;
    END
    ANTENNADIFFAREA 0.7227 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 0.6150 1.7700 0.7050 2.0800 ;
        RECT 1.9500 1.4450 2.1200 2.0800 ;
        RECT 2.4700 1.4450 2.6400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8750 1.8300 1.4850 1.9200 ;
      RECT 1.3950 1.4900 1.4850 1.8300 ;
      RECT 0.3550 1.4600 0.9650 1.5500 ;
      RECT 0.8750 1.5500 0.9650 1.8300 ;
      RECT 0.3550 1.5500 0.4450 1.8900 ;
      RECT 1.7050 0.4800 2.4000 0.5700 ;
      RECT 0.0950 0.7600 1.7950 0.8500 ;
      RECT 1.7050 0.5700 1.7950 0.7600 ;
      RECT 0.0950 0.4200 0.1850 0.7600 ;
      RECT 0.6150 0.4200 0.7050 0.7600 ;
      RECT 1.1350 0.4200 1.2250 0.7600 ;
  END
END OAI21_X3M_A12TH

MACRO OAI21_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7050 ;
        RECT 0.8750 0.3200 0.9650 0.7050 ;
        RECT 1.3950 0.3200 1.4850 0.7050 ;
        RECT 1.9150 0.3200 2.0050 0.7050 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3150 1.0500 0.9650 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3600 1.0500 2.0250 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3000 1.0500 2.9100 1.1500 ;
    END
    ANTENNAGATEAREA 0.2559 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9500 3.1500 1.2500 ;
        RECT 1.3900 1.2500 3.1500 1.3500 ;
        RECT 2.4350 0.8500 3.1500 0.9500 ;
        RECT 1.3950 1.3500 1.4850 1.7050 ;
        RECT 1.9150 1.3500 2.0050 1.7050 ;
        RECT 2.4300 1.3500 2.5200 1.7050 ;
        RECT 2.9550 1.3500 3.0450 1.7050 ;
        RECT 2.4350 0.6800 2.5250 0.8500 ;
        RECT 2.9550 0.6800 3.0450 0.8500 ;
    END
    ANTENNADIFFAREA 0.8286 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 2.6950 1.4950 2.7850 2.0800 ;
        RECT 3.2200 1.4950 3.3100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1350 1.8200 2.2650 1.9200 ;
      RECT 2.1750 1.4900 2.2650 1.8200 ;
      RECT 1.1350 1.3750 1.2250 1.8200 ;
      RECT 0.0950 1.2850 1.2250 1.3750 ;
      RECT 1.6550 1.4900 1.7450 1.8200 ;
      RECT 0.0950 1.3750 0.1850 1.7200 ;
      RECT 0.6150 1.3750 0.7050 1.7200 ;
      RECT 2.1750 0.4800 3.3050 0.5700 ;
      RECT 3.2150 0.5700 3.3050 0.6900 ;
      RECT 0.0950 0.7950 2.2650 0.8850 ;
      RECT 2.1750 0.5700 2.2650 0.7950 ;
      RECT 0.0950 0.4600 0.1850 0.7950 ;
      RECT 0.6150 0.4600 0.7050 0.7950 ;
      RECT 1.1350 0.4600 1.2250 0.7950 ;
      RECT 1.6550 0.4600 1.7450 0.7950 ;
  END
END OAI21_X4M_A12TH

MACRO OAI21_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.5600 ;
        RECT 0.8200 0.3200 0.9900 0.5600 ;
        RECT 1.3400 0.3200 1.5100 0.5600 ;
        RECT 1.8600 0.3200 2.0300 0.5600 ;
        RECT 2.3800 0.3200 2.5500 0.5600 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.2500 3.1350 1.3500 ;
        RECT 0.9850 1.1500 1.0850 1.2500 ;
        RECT 2.0250 1.1500 2.1250 1.2500 ;
        RECT 0.2350 1.0450 0.3250 1.2500 ;
        RECT 3.0450 1.0000 3.1350 1.2500 ;
        RECT 0.9850 1.0500 1.3750 1.1500 ;
        RECT 2.0250 1.0500 2.4050 1.1500 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5950 1.4500 4.3500 1.5500 ;
        RECT 0.5950 1.5500 0.6950 1.8800 ;
        RECT 1.6350 1.5500 1.7350 1.8800 ;
        RECT 2.6750 1.5500 2.7750 1.8800 ;
        RECT 3.6450 1.5500 3.7450 1.8800 ;
        RECT 4.1650 1.5500 4.2650 1.8800 ;
        RECT 4.2500 0.9600 4.3500 1.4500 ;
        RECT 4.2500 0.9500 4.5250 0.9600 ;
        RECT 3.3500 0.8500 4.5250 0.9500 ;
        RECT 3.3500 0.6600 3.5200 0.8500 ;
        RECT 3.8700 0.6600 4.0400 0.8500 ;
        RECT 4.4250 0.5300 4.5250 0.8500 ;
    END
    ANTENNADIFFAREA 1.2296 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4100 1.0500 4.1450 1.1800 ;
    END
    ANTENNAGATEAREA 0.3846 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0500 0.8350 1.1500 ;
        RECT 0.7450 0.9500 0.8350 1.0500 ;
        RECT 0.7450 0.8500 2.6050 0.9500 ;
        RECT 2.5150 0.9500 2.6050 1.0600 ;
        RECT 1.4850 0.9500 1.5850 1.0500 ;
        RECT 2.5150 1.0600 2.9050 1.1500 ;
        RECT 1.4850 1.0500 1.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.0750 1.7800 0.1750 2.0800 ;
        RECT 1.1150 1.7800 1.2150 2.0800 ;
        RECT 2.1550 1.7800 2.2550 2.0800 ;
        RECT 3.2750 1.7800 3.3750 2.0800 ;
        RECT 3.9050 1.6550 4.0050 2.0800 ;
        RECT 4.4250 1.6200 4.5250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.6750 0.4800 4.3200 0.5700 ;
      RECT 0.0750 0.6500 2.7750 0.7400 ;
      RECT 2.6750 0.5700 2.7750 0.6500 ;
      RECT 0.0750 0.5300 0.1750 0.6500 ;
      RECT 0.5600 0.4100 0.7300 0.6500 ;
      RECT 1.0800 0.4150 1.2500 0.6500 ;
      RECT 1.6000 0.4150 1.7700 0.6500 ;
      RECT 2.1200 0.4150 2.2900 0.6500 ;
  END
END OAI21_X6M_A12TH

MACRO OAI21_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4550 0.5800 ;
        RECT 0.8750 0.3200 0.9750 0.5800 ;
        RECT 1.3950 0.3200 1.4950 0.5800 ;
        RECT 1.9150 0.3200 2.0150 0.5800 ;
        RECT 2.4350 0.3200 2.5350 0.5800 ;
        RECT 2.9550 0.3200 3.0550 0.5800 ;
        RECT 3.4750 0.3200 3.5750 0.5800 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.0500 0.8550 1.1500 ;
        RECT 0.7650 0.9500 0.8550 1.0500 ;
        RECT 0.7650 0.8500 3.6650 0.9500 ;
        RECT 1.5150 0.9500 1.6150 1.0500 ;
        RECT 2.5550 0.9500 2.6550 1.0500 ;
        RECT 3.5750 0.9500 3.6650 1.0500 ;
        RECT 1.5150 1.0500 1.8850 1.1500 ;
        RECT 2.5550 1.0500 2.9250 1.1500 ;
        RECT 3.5750 1.0500 3.9650 1.1500 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4950 1.0500 5.7750 1.1500 ;
    END
    ANTENNAGATEAREA 0.5115 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.2500 4.1950 1.3500 ;
        RECT 1.0050 1.1500 1.1050 1.2500 ;
        RECT 2.0350 1.1500 2.1350 1.2500 ;
        RECT 3.0750 1.1500 3.1750 1.2500 ;
        RECT 4.1050 1.0500 4.1950 1.2500 ;
        RECT 0.2550 1.0450 0.3450 1.2500 ;
        RECT 1.0050 1.0500 1.3750 1.1500 ;
        RECT 2.0350 1.0500 2.4050 1.1500 ;
        RECT 3.0750 1.0500 3.4450 1.1500 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 1.4500 6.1500 1.5800 ;
        RECT 0.6150 1.5800 0.7150 1.8800 ;
        RECT 1.6550 1.5800 1.7550 1.8850 ;
        RECT 2.6950 1.5800 2.7950 1.8800 ;
        RECT 3.7350 1.5800 3.8350 1.8800 ;
        RECT 4.9550 1.5800 5.0550 1.8600 ;
        RECT 5.4750 1.5800 5.5750 1.8800 ;
        RECT 5.9950 1.5800 6.1500 1.8800 ;
        RECT 6.0000 0.6100 6.1500 1.4500 ;
        RECT 4.3800 0.4800 6.1500 0.6100 ;
    END
    ANTENNADIFFAREA 1.6953 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.0950 1.7700 0.1950 2.0800 ;
        RECT 1.1350 1.7700 1.2350 2.0800 ;
        RECT 2.1750 1.7700 2.2750 2.0800 ;
        RECT 3.2150 1.7700 3.3150 2.0800 ;
        RECT 4.4900 1.7700 4.5900 2.0800 ;
        RECT 5.2150 1.6700 5.3150 2.0800 ;
        RECT 5.7350 1.6700 5.8350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.1750 0.7900 5.8900 0.8800 ;
      RECT 4.1750 0.7600 4.2750 0.7900 ;
      RECT 0.1000 0.6700 4.2750 0.7600 ;
      RECT 4.1750 0.4500 4.2750 0.6700 ;
      RECT 3.7400 0.4100 3.8300 0.6700 ;
      RECT 0.1000 0.5500 0.1900 0.6700 ;
      RECT 0.6200 0.4100 0.7100 0.6700 ;
      RECT 1.1400 0.4100 1.2300 0.6700 ;
      RECT 1.6600 0.4100 1.7500 0.6700 ;
      RECT 2.1800 0.4100 2.2700 0.6700 ;
      RECT 2.7000 0.4100 2.7900 0.6700 ;
      RECT 3.2200 0.4100 3.3100 0.6700 ;
  END
END OAI21_X8M_A12TH

MACRO OAI221_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6900 ;
        RECT 0.6350 0.3200 0.8050 0.3950 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5100 1.6500 1.7500 1.7500 ;
        RECT 1.5900 1.7500 1.7500 1.7550 ;
        RECT 0.5100 1.7500 0.6800 1.9400 ;
        RECT 0.7900 1.7500 0.9600 1.9900 ;
        RECT 1.6500 0.9600 1.7500 1.6500 ;
        RECT 1.5900 1.7550 1.6800 1.8750 ;
        RECT 1.5900 0.8700 1.7500 0.9600 ;
        RECT 1.5900 0.5900 1.6800 0.8700 ;
    END
    ANTENNADIFFAREA 0.24935 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.0500 1.5250 1.1500 ;
        RECT 1.4350 1.1500 1.5250 1.2700 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END C0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0000 1.2500 1.2950 1.3500 ;
        RECT 1.2050 1.3500 1.2950 1.4900 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7100 1.4500 1.0350 1.5500 ;
        RECT 0.8000 1.3400 0.8900 1.4500 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3700 1.2500 0.6900 1.3500 ;
        RECT 0.4450 1.3500 0.5350 1.4650 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8100 0.3700 1.1400 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.2650 1.8400 1.4350 2.0800 ;
        RECT 0.0800 1.6300 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6100 1.0200 1.1000 1.1100 ;
      RECT 1.0100 0.9550 1.1000 1.0200 ;
      RECT 0.6100 0.7000 0.7000 1.0200 ;
      RECT 1.0100 0.6650 1.2000 0.9550 ;
      RECT 0.3000 0.6100 0.7000 0.7000 ;
      RECT 0.3000 0.4100 0.4700 0.6100 ;
      RECT 0.8100 0.5750 0.9000 0.9300 ;
      RECT 0.8100 0.4850 1.4200 0.5750 ;
      RECT 1.3300 0.5750 1.4200 0.9300 ;
  END
END OAI221_X0P5M_A12TH

MACRO OAI221_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7850 ;
        RECT 0.6000 0.3200 0.6900 0.7850 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9800 0.1650 1.1000 ;
        RECT 0.0500 1.1000 0.2750 1.1900 ;
        RECT 0.1850 1.1900 0.2750 1.3100 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3650 1.2500 0.6300 1.3500 ;
        RECT 0.4250 1.0650 0.5150 1.2500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2600 1.0950 1.3900 ;
        RECT 1.0050 1.3900 1.0950 1.4700 ;
        RECT 0.8500 1.1950 0.9800 1.2600 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.4500 1.4950 1.5500 ;
        RECT 1.2350 1.2800 1.3250 1.4500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END B1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 0.9600 1.5550 1.3400 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.6500 1.7500 1.7500 ;
        RECT 0.4900 1.7500 0.6600 1.9550 ;
        RECT 0.8600 1.7500 1.0300 1.9550 ;
        RECT 1.6200 1.7500 1.7100 1.8600 ;
        RECT 1.6500 0.8400 1.7500 1.6500 ;
        RECT 1.6300 0.7800 1.7500 0.8400 ;
        RECT 1.6300 0.4700 1.7200 0.7800 ;
    END
    ANTENNADIFFAREA 0.3885 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.3100 1.8600 1.4800 2.0800 ;
        RECT 0.0800 1.6600 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.8750 1.2400 0.9650 ;
      RECT 1.0700 0.6650 1.2400 0.8750 ;
      RECT 0.3400 0.5950 0.4300 0.8750 ;
      RECT 0.8500 0.5750 0.9400 0.7850 ;
      RECT 0.8500 0.4850 1.4600 0.5750 ;
      RECT 1.3700 0.5750 1.4600 0.8550 ;
      RECT 0.8500 0.4150 0.9400 0.4850 ;
  END
END OAI221_X0P7M_A12TH

MACRO OAI221_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6300 ;
        RECT 0.6000 0.3200 0.6900 0.6300 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.0500 1.1100 1.1500 ;
        RECT 0.7900 1.1500 0.8800 1.2700 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.2950 1.2050 ;
        RECT 0.2050 1.2050 0.2950 1.2600 ;
        RECT 0.0500 1.0100 0.1500 1.0500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3850 1.2500 0.6250 1.3700 ;
        RECT 0.4450 1.0700 0.5450 1.2500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9900 1.2500 1.3200 1.3400 ;
        RECT 0.9900 1.3400 1.2300 1.3500 ;
        RECT 1.2300 1.0500 1.3200 1.2500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END B1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0000 1.5500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9000 1.7500 1.5300 ;
        RECT 0.5550 1.5300 1.7500 1.6300 ;
        RECT 1.6300 0.8400 1.7500 0.9000 ;
        RECT 1.6050 1.6300 1.7500 1.7100 ;
        RECT 0.5550 1.6300 0.6550 1.9000 ;
        RECT 0.8800 1.6300 0.9800 1.9000 ;
        RECT 1.6300 0.4700 1.7200 0.8400 ;
        RECT 1.6050 1.7100 1.6950 1.9900 ;
    END
    ANTENNADIFFAREA 0.4962 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.1000 1.7700 0.1900 2.0800 ;
        RECT 1.3450 1.7200 1.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.8700 1.2400 0.9600 ;
      RECT 1.0700 0.6650 1.2400 0.8700 ;
      RECT 0.3400 0.5900 0.4300 0.8700 ;
      RECT 0.8500 0.5700 0.9400 0.7800 ;
      RECT 0.8500 0.4800 1.4600 0.5700 ;
      RECT 1.3700 0.5700 1.4600 0.8500 ;
      RECT 0.8500 0.4100 0.9400 0.4800 ;
  END
END OAI221_X1M_A12TH

MACRO OAI221_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.6850 ;
        RECT 0.8350 0.3200 1.0050 0.6850 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4900 1.0500 1.9100 1.1500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 1.1650 1.3500 ;
        RECT 0.2500 1.1350 0.3400 1.2500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.0500 0.9100 1.1500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2900 1.2500 2.2200 1.3500 ;
        RECT 1.2900 1.1200 1.3800 1.2500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END B1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3400 1.0500 2.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 1.4500 3.1150 1.5500 ;
        RECT 0.6150 1.5500 0.7050 1.9800 ;
        RECT 1.6550 1.5500 1.7450 1.9800 ;
        RECT 2.4250 1.5500 2.5950 1.9000 ;
        RECT 2.9450 1.5500 3.1150 1.9000 ;
        RECT 2.8500 0.8550 2.9500 1.4500 ;
        RECT 2.6650 0.7550 2.9500 0.8550 ;
    END
    ANTENNADIFFAREA 0.4746 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0950 1.7350 0.1850 2.0800 ;
        RECT 1.1350 1.7350 1.2250 2.0800 ;
        RECT 2.1750 1.7350 2.2650 2.0800 ;
        RECT 2.7250 1.6700 2.8150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.4650 0.4800 3.1350 0.5700 ;
      RECT 1.3950 0.8600 2.5550 0.9500 ;
      RECT 1.3950 0.7000 1.4850 0.8600 ;
      RECT 1.9150 0.7000 2.0050 0.8600 ;
      RECT 2.4650 0.5700 2.5550 0.8600 ;
      RECT 0.0950 0.8000 1.2250 0.8900 ;
      RECT 1.1350 0.5700 1.2250 0.8000 ;
      RECT 1.1350 0.4800 2.3050 0.5700 ;
      RECT 1.6150 0.5700 1.7850 0.7700 ;
      RECT 2.1350 0.5700 2.3050 0.7700 ;
      RECT 0.0950 0.4400 0.1850 0.8000 ;
      RECT 0.6150 0.4400 0.7050 0.8000 ;
  END
END OAI221_X1P4M_A12TH

MACRO OAI221_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6400 ;
        RECT 0.8750 0.3200 0.9650 0.6400 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5200 1.0500 1.9450 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.2500 1.1250 1.3500 ;
        RECT 0.1950 1.0500 0.2950 1.2500 ;
        RECT 1.0250 1.0500 1.1250 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5100 1.0500 2.9300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.8750 3.1500 1.4500 ;
        RECT 0.6150 1.4500 3.1500 1.5500 ;
        RECT 2.6700 0.7750 3.1500 0.8750 ;
        RECT 0.6150 1.5500 0.7050 1.8800 ;
        RECT 1.6550 1.5500 1.7450 1.8800 ;
        RECT 2.4650 1.5500 2.5550 1.8800 ;
        RECT 2.9850 1.5500 3.0750 1.8800 ;
    END
    ANTENNADIFFAREA 0.6555 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 2.1750 1.7700 2.2650 2.0800 ;
        RECT 2.7250 1.7100 2.8150 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2850 1.2500 2.1900 1.3500 ;
        RECT 1.2850 1.0500 1.3850 1.2500 ;
        RECT 2.1000 1.0500 2.1900 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END B1
  OBS
    LAYER M1 ;
      RECT 0.0950 0.8300 1.2250 0.9200 ;
      RECT 1.1350 0.5700 1.2250 0.8300 ;
      RECT 1.1350 0.4800 2.3050 0.5700 ;
      RECT 1.6150 0.5700 1.7850 0.7700 ;
      RECT 2.1350 0.5700 2.3050 0.7700 ;
      RECT 0.0950 0.4800 0.1850 0.8300 ;
      RECT 0.6150 0.4800 0.7050 0.8300 ;
      RECT 2.4650 0.4800 3.1400 0.5700 ;
      RECT 1.3950 0.8600 2.5550 0.9500 ;
      RECT 1.3950 0.7400 1.4850 0.8600 ;
      RECT 1.9150 0.7400 2.0050 0.8600 ;
      RECT 2.4650 0.5700 2.5550 0.8600 ;
  END
END OAI221_X2M_A12TH

MACRO OAI221_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6300 ;
        RECT 0.8750 0.3200 0.9650 0.6300 ;
        RECT 1.3950 0.3200 1.4850 0.6300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1350 1.2500 4.3800 1.3500 ;
        RECT 1.1350 1.3500 1.2250 1.7300 ;
        RECT 1.6550 1.3500 1.7450 1.7300 ;
        RECT 2.1750 1.3500 2.2650 1.7300 ;
        RECT 3.5500 1.3500 3.6400 1.7700 ;
        RECT 4.0700 1.3500 4.1600 1.7700 ;
        RECT 4.2800 0.5800 4.3800 1.2500 ;
        RECT 3.7250 0.4800 4.3800 0.5800 ;
        RECT 3.7250 0.5800 3.8950 0.7700 ;
    END
    ANTENNADIFFAREA 0.9735 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4400 1.0500 3.9300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END C0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.0500 3.1600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8400 1.0500 2.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.0500 1.5600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0500 0.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 0.6150 1.7700 0.7050 2.0800 ;
        RECT 2.6950 1.7700 2.7850 2.0800 ;
        RECT 3.2150 1.7700 3.3050 2.0800 ;
        RECT 3.7700 1.4700 3.9400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8750 1.8300 1.4850 1.9200 ;
      RECT 1.3950 1.4850 1.4850 1.8300 ;
      RECT 0.8750 1.4300 0.9650 1.8300 ;
      RECT 0.3550 1.3400 0.9650 1.4300 ;
      RECT 0.3550 1.4300 0.4450 1.7700 ;
      RECT 2.4350 1.4900 3.0450 1.5800 ;
      RECT 2.9550 1.5800 3.0450 1.9200 ;
      RECT 1.9150 1.8300 2.5250 1.9200 ;
      RECT 2.4350 1.5800 2.5250 1.8300 ;
      RECT 1.9150 1.4850 2.0050 1.8300 ;
      RECT 0.0950 0.8300 1.7450 0.9200 ;
      RECT 1.6550 0.5700 1.7450 0.8300 ;
      RECT 1.6550 0.4800 3.3450 0.5700 ;
      RECT 2.1350 0.5700 2.3050 0.7700 ;
      RECT 2.6550 0.5700 2.8250 0.7700 ;
      RECT 3.1750 0.5700 3.3450 0.7700 ;
      RECT 0.0950 0.4850 0.1850 0.8300 ;
      RECT 0.6150 0.4850 0.7050 0.8300 ;
      RECT 1.1350 0.4850 1.2250 0.8300 ;
      RECT 1.9150 0.8650 4.1150 0.9550 ;
      RECT 4.0250 0.7450 4.1150 0.8650 ;
      RECT 1.9150 0.7450 2.0050 0.8650 ;
      RECT 2.4350 0.7450 2.5250 0.8650 ;
      RECT 2.9550 0.7450 3.0450 0.8650 ;
      RECT 3.5050 0.5250 3.5950 0.8650 ;
  END
END OAI221_X3M_A12TH

MACRO OAI221_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6300 ;
        RECT 0.6150 0.3200 0.7050 0.6300 ;
        RECT 1.1350 0.3200 1.2250 0.6300 ;
        RECT 1.6550 0.3200 1.7450 0.6300 ;
        RECT 2.1750 0.3200 2.2650 0.6300 ;
    END
  END VSS

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7300 1.0500 5.2200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 0.8100 5.5500 1.4500 ;
        RECT 0.6150 1.4500 5.5500 1.5500 ;
        RECT 4.7550 0.7100 5.5500 0.8100 ;
        RECT 0.6150 1.5500 0.7050 1.8800 ;
        RECT 1.6550 1.5500 1.7450 1.8800 ;
        RECT 2.9850 1.5500 3.0750 1.8800 ;
        RECT 4.0250 1.5500 4.1150 1.8800 ;
        RECT 4.8800 1.5500 4.9700 1.8800 ;
        RECT 5.4000 1.5500 5.4900 1.8800 ;
    END
    ANTENNADIFFAREA 1.239 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.2500 4.5350 1.3500 ;
        RECT 3.3900 1.1600 3.7600 1.2500 ;
        RECT 2.6400 1.0500 2.7400 1.2500 ;
        RECT 4.4350 1.0500 4.5350 1.2500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.2500 2.1700 1.3500 ;
        RECT 1.0200 1.1600 1.3900 1.2500 ;
        RECT 0.2550 1.0500 0.3550 1.2500 ;
        RECT 2.0700 1.0500 2.1700 1.2500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.0500 0.8900 1.1500 ;
        RECT 0.7900 1.0400 0.8900 1.0500 ;
        RECT 0.7900 0.9400 1.6200 1.0400 ;
        RECT 1.5200 1.0400 1.6200 1.0500 ;
        RECT 1.5200 1.0500 1.9300 1.1500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 2.1800 1.7700 2.2700 2.0800 ;
        RECT 2.4650 1.7700 2.5550 2.0800 ;
        RECT 3.5050 1.7700 3.5950 2.0800 ;
        RECT 4.5450 1.7700 4.6350 2.0800 ;
        RECT 5.1400 1.7300 5.2300 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0500 3.2550 1.1500 ;
        RECT 3.1550 1.0400 3.2550 1.0500 ;
        RECT 3.1550 0.9400 3.9850 1.0400 ;
        RECT 3.8850 1.0400 3.9850 1.0500 ;
        RECT 3.8850 1.0500 4.2950 1.1500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.3550 0.7500 4.4250 0.8400 ;
      RECT 0.3550 0.4100 0.4450 0.7500 ;
      RECT 0.8750 0.4100 0.9650 0.7500 ;
      RECT 1.3950 0.4100 1.4850 0.7500 ;
      RECT 1.9150 0.4100 2.0050 0.7500 ;
      RECT 2.4050 0.4800 5.7300 0.5700 ;
      RECT 4.5450 0.5700 4.6350 0.9100 ;
  END
END OAI221_X4M_A12TH

MACRO OAI222_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 1.3100 0.3200 1.4000 0.5050 ;
        RECT 1.8300 0.3200 1.9200 0.5800 ;
    END
  END VSS

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END C0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5200 1.0500 0.8450 1.1500 ;
        RECT 0.5200 1.1500 0.6100 1.2700 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END C1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9650 1.0500 1.2750 1.1500 ;
        RECT 1.1850 1.1500 1.2750 1.2800 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0500 1.5500 1.4700 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8400 0.8500 1.9500 1.2400 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.6500 1.4550 1.7500 ;
        RECT 0.0800 1.7500 0.1700 1.9900 ;
        RECT 1.1250 1.7500 1.2150 1.9900 ;
        RECT 1.3650 1.5600 1.4550 1.6500 ;
        RECT 0.3400 0.6600 0.4300 1.6500 ;
    END
    ANTENNADIFFAREA 0.289625 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.5650 1.8400 0.7350 2.0800 ;
        RECT 1.8300 1.3600 1.9200 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7100 1.2500 1.0950 1.3600 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END B1
  OBS
    LAYER M1 ;
      RECT 0.0800 0.4800 1.2150 0.5700 ;
      RECT 0.6050 0.5700 0.6950 0.9300 ;
      RECT 1.1250 0.5700 1.2150 0.7800 ;
      RECT 0.0800 0.5700 0.1700 0.9450 ;
      RECT 0.8650 0.8700 1.6600 0.9600 ;
      RECT 1.5700 0.4100 1.6600 0.8700 ;
      RECT 0.8650 0.6600 0.9550 0.8700 ;
  END
END OAI222_X0P5M_A12TH

MACRO OAI222_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.7200 ;
    END
  END VSS

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7800 0.9950 1.9500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END C1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0100 0.5550 1.3950 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9750 1.5600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END C0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.0300 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6900 1.0500 1.1100 1.1500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.8800 2.1500 1.4500 ;
        RECT 0.6300 1.4500 2.1500 1.5500 ;
        RECT 1.7000 0.7800 2.1500 0.8800 ;
        RECT 0.6300 1.5500 0.7300 1.8650 ;
        RECT 1.4400 1.5500 1.5400 1.8650 ;
        RECT 1.7000 0.6700 1.8000 0.7800 ;
    END
    ANTENNADIFFAREA 0.3469 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8950 1.2500 1.3150 1.3500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.1050 1.6550 0.1950 2.0800 ;
        RECT 1.1600 1.6550 1.2500 2.0800 ;
        RECT 1.8950 1.6550 1.9850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1050 0.8100 1.2500 0.9000 ;
      RECT 1.1600 0.6750 1.2500 0.8100 ;
      RECT 0.6350 0.4750 0.7250 0.8100 ;
      RECT 0.1050 0.4750 0.1950 0.8100 ;
      RECT 0.9000 0.4800 2.0550 0.5700 ;
      RECT 1.9650 0.5700 2.0550 0.6900 ;
      RECT 0.9000 0.5700 0.9900 0.6900 ;
      RECT 1.4450 0.5700 1.5350 0.8850 ;
  END
END OAI222_X0P7M_A12TH

MACRO OAI222_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.6300 ;
    END
  END VSS

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0600 1.1900 1.4000 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.7600 2.1500 1.5650 ;
        RECT 0.6300 1.5650 2.1500 1.6650 ;
        RECT 1.6450 0.6600 2.1500 0.7600 ;
        RECT 0.6300 1.6650 0.7300 1.9750 ;
        RECT 1.4400 1.6650 1.5400 1.9900 ;
    END
    ANTENNADIFFAREA 0.4894 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0100 0.8100 1.3100 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1600 1.5550 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0100 1.5900 1.3650 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END C0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0750 0.5500 1.5150 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8450 0.8900 1.9550 1.3300 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END C1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.1050 1.7700 0.1950 2.0800 ;
        RECT 1.1600 1.7700 1.2500 2.0800 ;
        RECT 1.9650 1.7700 2.0550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1050 0.7700 1.3100 0.8600 ;
      RECT 0.6350 0.4300 0.7250 0.7700 ;
      RECT 0.1050 0.4300 0.1950 0.7700 ;
      RECT 0.8400 0.4800 2.1050 0.5700 ;
      RECT 1.4450 0.5700 1.5350 0.8900 ;
  END
END OAI222_X1M_A12TH

MACRO OAI222_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6000 ;
        RECT 0.6000 0.3200 0.6900 0.6000 ;
        RECT 1.1200 0.3200 1.2100 0.5450 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.4500 1.0550 1.5500 ;
        RECT 0.2350 1.3200 0.3250 1.4500 ;
        RECT 0.9650 1.3200 1.0550 1.4500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4350 1.0500 0.8550 1.1500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.4500 2.3000 1.5500 ;
        RECT 1.4100 1.3200 1.5000 1.4500 ;
        RECT 2.2100 1.3200 2.3000 1.4500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6100 1.2500 2.0950 1.3500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END B0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5700 1.4500 3.4150 1.5500 ;
        RECT 2.5700 1.3200 2.6600 1.4500 ;
        RECT 3.3250 1.3200 3.4150 1.4500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END C1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7700 1.2500 3.1900 1.3500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.6500 3.0400 1.7500 ;
        RECT 0.5600 1.7500 0.7300 1.9400 ;
        RECT 1.8300 1.7500 2.0000 1.9400 ;
        RECT 2.8700 1.7500 3.0400 1.9400 ;
        RECT 2.3900 1.0450 2.4800 1.6500 ;
        RECT 2.3900 0.9550 3.2200 1.0450 ;
        RECT 2.6100 0.6650 2.7800 0.9550 ;
        RECT 3.1300 0.6650 3.3000 0.9550 ;
    END
    ANTENNADIFFAREA 0.584 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 1.0200 1.8800 1.1900 2.0800 ;
        RECT 1.3700 1.8800 1.5400 2.0800 ;
        RECT 2.3500 1.8800 2.5200 2.0800 ;
        RECT 0.1350 1.8400 0.2350 2.0800 ;
        RECT 3.3650 1.8400 3.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1100 1.0250 2.1800 1.1150 ;
      RECT 2.0900 0.9550 2.1800 1.0250 ;
      RECT 1.1100 0.8000 1.2000 1.0250 ;
      RECT 1.5700 0.6650 1.7400 1.0250 ;
      RECT 2.0900 0.6650 2.2600 0.9550 ;
      RECT 0.3000 0.7000 1.2000 0.8000 ;
      RECT 0.3000 0.4400 0.4700 0.7000 ;
      RECT 0.8200 0.4400 0.9900 0.7000 ;
      RECT 1.3900 0.4850 3.5200 0.5750 ;
      RECT 3.4300 0.5750 3.5200 0.8550 ;
      RECT 1.3100 0.6450 1.4800 0.9350 ;
      RECT 1.3900 0.5750 1.4800 0.6450 ;
      RECT 1.8700 0.5750 1.9600 0.8550 ;
      RECT 2.3900 0.5750 2.4800 0.8550 ;
      RECT 2.9100 0.5750 3.0000 0.8550 ;
  END
END OAI222_X1P4M_A12TH

MACRO OAI222_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6400 ;
        RECT 0.8750 0.3200 0.9650 0.6200 ;
    END
  END VSS

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.2900 3.5600 1.3900 ;
        RECT 2.6500 1.0400 2.7500 1.2900 ;
        RECT 3.4600 1.0400 3.5600 1.2900 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END C1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0100 1.3850 1.2500 ;
        RECT 1.2500 1.2500 2.2000 1.3500 ;
        RECT 2.1000 1.0550 2.2000 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5400 1.0500 1.9600 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8800 1.0500 3.3100 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END C0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.2500 1.1500 1.3500 ;
        RECT 0.1950 1.0550 0.2950 1.2500 ;
        RECT 1.0500 1.0550 1.1500 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.4500 2.5500 1.5500 ;
        RECT 2.4500 1.5500 3.0900 1.6500 ;
        RECT 0.6100 1.5500 0.7100 1.8800 ;
        RECT 1.6500 1.5500 1.7500 1.8800 ;
        RECT 2.4500 0.8300 2.5500 1.4500 ;
        RECT 2.9900 1.6500 3.0900 1.9600 ;
        RECT 2.4500 0.7300 3.4050 0.8300 ;
    END
    ANTENNADIFFAREA 0.824 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.0950 1.7650 0.1850 2.0800 ;
        RECT 2.1750 1.7650 2.2650 2.0800 ;
        RECT 2.4750 1.7650 2.5650 2.0800 ;
        RECT 3.5150 1.7650 3.6050 2.0800 ;
        RECT 1.1350 1.7600 1.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 0.7350 2.3250 0.8250 ;
      RECT 1.1350 0.4150 1.2250 0.7350 ;
      RECT 0.0950 0.4150 0.1850 0.7350 ;
      RECT 0.6150 0.4150 0.7050 0.7350 ;
      RECT 3.5150 0.5700 3.6050 0.8900 ;
      RECT 1.3350 0.4800 3.6050 0.5700 ;
  END
END OAI222_X2M_A12TH

MACRO OAI222_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6100 ;
        RECT 0.8750 0.3200 0.9650 0.6100 ;
        RECT 1.3950 0.3200 1.4850 0.6100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 1.1350 1.7850 1.2250 2.0800 ;
        RECT 2.1750 1.7850 2.2650 2.0800 ;
        RECT 3.2150 1.7850 3.3050 2.0800 ;
        RECT 4.0150 1.7850 4.1050 2.0800 ;
        RECT 0.0950 1.7650 0.1850 2.0800 ;
        RECT 5.0550 1.7650 5.1450 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.0100 0.3550 1.2900 ;
        RECT 0.2250 1.2900 1.0500 1.3900 ;
        RECT 0.9500 1.2300 1.0500 1.2900 ;
        RECT 0.9500 1.1300 1.3600 1.2300 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0100 1.5800 1.2650 ;
        RECT 0.7500 0.9100 1.5800 1.0100 ;
        RECT 0.7500 1.0100 0.8500 1.0550 ;
        RECT 0.4500 1.0550 0.8500 1.1550 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 1.0350 3.1500 1.2650 ;
        RECT 2.2400 0.9350 3.1500 1.0350 ;
        RECT 2.2400 1.0350 2.3400 1.0850 ;
        RECT 1.9700 1.0850 2.3400 1.1850 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END B1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 1.0100 3.7500 1.2900 ;
        RECT 3.6500 1.2900 4.4500 1.3900 ;
        RECT 4.3500 1.2300 4.4500 1.2900 ;
        RECT 4.3500 1.1300 4.7600 1.2300 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END C0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.0450 5.0000 1.2650 ;
        RECT 4.8500 0.9900 4.9500 1.0450 ;
        RECT 4.1600 0.8900 4.9500 0.9900 ;
        RECT 4.1600 0.9900 4.2600 1.0500 ;
        RECT 3.8500 1.0500 4.2600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.8000 3.5500 1.5750 ;
        RECT 0.6100 1.5750 4.6300 1.6750 ;
        RECT 3.4500 0.7000 4.9450 0.8000 ;
        RECT 0.6100 1.6750 0.7100 1.9900 ;
        RECT 1.6500 1.6750 1.7500 1.9900 ;
        RECT 2.6900 1.6750 2.7900 1.9900 ;
        RECT 3.4900 1.6750 3.5900 1.9900 ;
        RECT 4.5300 1.6750 4.6300 1.9900 ;
    END
    ANTENNADIFFAREA 1.3005 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7550 1.2900 2.5500 1.3900 ;
        RECT 2.4500 1.2350 2.5500 1.2900 ;
        RECT 1.7550 1.0100 1.8550 1.2900 ;
        RECT 2.4500 1.1350 2.9200 1.2350 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.0950 0.7300 3.3600 0.8200 ;
      RECT 1.6550 0.4100 1.7450 0.7300 ;
      RECT 0.0950 0.4100 0.1850 0.7300 ;
      RECT 0.6150 0.4100 0.7050 0.7300 ;
      RECT 1.1350 0.4100 1.2250 0.7300 ;
      RECT 5.0550 0.5700 5.1450 0.9000 ;
      RECT 1.8550 0.4800 5.1450 0.5700 ;
  END
END OAI222_X3M_A12TH

MACRO OAI222_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6300 ;
        RECT 0.8750 0.3200 0.9650 0.6300 ;
        RECT 1.3950 0.3200 1.4850 0.6300 ;
        RECT 1.9150 0.3200 2.0050 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 2.1750 1.7700 2.2650 2.0800 ;
        RECT 3.2150 1.7700 3.3050 2.0800 ;
        RECT 4.2550 1.7700 4.3450 2.0800 ;
        RECT 4.5350 1.7700 4.6250 2.0800 ;
        RECT 5.5750 1.7700 5.6650 2.0800 ;
        RECT 6.6150 1.7700 6.7050 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.0500 0.8400 1.1500 ;
        RECT 0.7400 1.0250 0.8400 1.0500 ;
        RECT 0.7400 0.9250 1.5750 1.0250 ;
        RECT 1.4750 1.0250 1.5750 1.0500 ;
        RECT 1.4750 1.0500 1.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.2500 ;
        RECT 0.2500 1.2500 1.0500 1.3500 ;
        RECT 0.9500 1.2350 1.0500 1.2500 ;
        RECT 0.9500 1.1350 1.3600 1.2350 ;
        RECT 1.2600 1.2350 1.3600 1.2500 ;
        RECT 1.2600 1.2500 2.1150 1.3500 ;
        RECT 2.0150 1.0500 2.1150 1.2500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5100 1.0500 2.9150 1.1500 ;
        RECT 2.8150 1.0150 2.9150 1.0500 ;
        RECT 2.8150 0.9150 3.6550 1.0150 ;
        RECT 3.5550 1.0150 3.6550 1.0500 ;
        RECT 3.5550 1.0500 3.9600 1.1500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0000 1.0500 5.2750 1.1500 ;
        RECT 5.1750 1.0200 5.2750 1.0500 ;
        RECT 5.1750 0.9200 6.0150 1.0200 ;
        RECT 5.9150 1.0200 6.0150 1.0500 ;
        RECT 5.9150 1.0500 6.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.8000 4.5500 1.4500 ;
        RECT 0.6100 1.4500 6.1900 1.5500 ;
        RECT 4.4500 0.7000 6.5050 0.8000 ;
        RECT 0.6100 1.5500 0.7100 1.8850 ;
        RECT 1.6500 1.5500 1.7500 1.8850 ;
        RECT 2.6900 1.5500 2.7900 1.8850 ;
        RECT 3.7300 1.5500 3.8300 1.8850 ;
        RECT 5.0500 1.5500 5.1500 1.8850 ;
        RECT 6.0900 1.5500 6.1900 1.8850 ;
    END
    ANTENNADIFFAREA 1.648 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.0100 2.3700 1.2500 ;
        RECT 2.2500 1.2500 3.1250 1.3500 ;
        RECT 3.0250 1.2250 3.1250 1.2500 ;
        RECT 3.0250 1.1350 3.4400 1.2250 ;
        RECT 3.3400 1.2250 3.4400 1.2500 ;
        RECT 3.3400 1.2500 4.1950 1.3500 ;
        RECT 4.0950 1.0500 4.1950 1.2500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.0100 4.7800 1.2500 ;
        RECT 4.6500 1.2500 5.4850 1.3500 ;
        RECT 5.3850 1.2250 5.4850 1.2500 ;
        RECT 5.3850 1.1350 5.8050 1.2250 ;
        RECT 5.7050 1.2250 5.8050 1.2550 ;
        RECT 5.7050 1.2550 6.5500 1.3450 ;
        RECT 6.4600 1.0500 6.5500 1.2550 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END C1
  OBS
    LAYER M1 ;
      RECT 4.2550 0.8200 4.3450 0.9400 ;
      RECT 0.0950 0.7300 4.3450 0.8200 ;
      RECT 0.0950 0.4100 0.1850 0.7300 ;
      RECT 0.6150 0.4100 0.7050 0.7300 ;
      RECT 1.1350 0.4100 1.2250 0.7300 ;
      RECT 1.6550 0.4100 1.7450 0.7300 ;
      RECT 6.6150 0.5700 6.7050 0.8900 ;
      RECT 2.3750 0.4800 6.7050 0.5700 ;
  END
END OAI222_X4M_A12TH

MACRO OAI22_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.9300 0.3200 1.0300 0.6800 ;
    END
  END VSS

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0100 0.9500 1.4300 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5750 1.4300 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 0.9800 1.3500 1.4000 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9000 0.3500 1.5900 ;
        RECT 0.2500 1.5900 0.7600 1.6900 ;
        RECT 0.2500 0.8000 0.5050 0.9000 ;
        RECT 0.6700 1.6900 0.7600 1.9600 ;
        RECT 0.4050 0.6600 0.5050 0.8000 ;
    END
    ANTENNADIFFAREA 0.152275 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1450 1.8000 0.2450 2.0800 ;
        RECT 1.1900 1.5750 1.2900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6750 0.7700 1.2850 0.8600 ;
      RECT 1.1950 0.6000 1.2850 0.7700 ;
      RECT 0.6750 0.5700 0.7650 0.7700 ;
      RECT 0.1500 0.4800 0.7650 0.5700 ;
      RECT 0.1500 0.5700 0.2400 0.7100 ;
  END
END OAI22_X0P5M_A12TH

MACRO OAI22_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.9350 0.3200 1.0250 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1500 1.6600 0.2400 2.0800 ;
        RECT 1.1950 1.6400 1.2850 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9000 0.3500 1.4500 ;
        RECT 0.2500 1.4500 0.7650 1.5500 ;
        RECT 0.2500 0.8000 0.5050 0.9000 ;
        RECT 0.6650 1.5500 0.7650 1.8800 ;
        RECT 0.4050 0.6650 0.5050 0.8000 ;
    END
    ANTENNADIFFAREA 0.216225 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 1.0000 1.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9700 0.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END B1
  OBS
    LAYER M1 ;
      RECT 0.6750 0.7700 1.2850 0.8600 ;
      RECT 1.1950 0.4650 1.2850 0.7700 ;
      RECT 0.6750 0.5750 0.7650 0.7700 ;
      RECT 0.1500 0.4850 0.7650 0.5750 ;
      RECT 0.1500 0.5750 0.2400 0.7100 ;
  END
END OAI22_X0P7M_A12TH

MACRO OAI22_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.5250 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9800 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.8800 0.5500 1.3150 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9900 0.7900 1.3900 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9800 1.1500 1.4000 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8700 1.3500 1.5800 ;
        RECT 0.6100 1.5800 1.3500 1.6800 ;
        RECT 0.8700 0.7700 1.3500 0.8700 ;
        RECT 0.6100 1.6800 0.7100 1.9900 ;
        RECT 0.8700 0.6600 0.9700 0.7700 ;
    END
    ANTENNADIFFAREA 0.30295 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0950 1.7900 0.1850 2.0800 ;
        RECT 1.1400 1.7900 1.2300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6150 0.4800 1.2400 0.5700 ;
      RECT 1.1500 0.5700 1.2400 0.6800 ;
      RECT 0.0950 0.6200 0.7050 0.7100 ;
      RECT 0.6150 0.5700 0.7050 0.6200 ;
      RECT 0.0950 0.7100 0.1850 0.8600 ;
      RECT 0.0950 0.4500 0.1850 0.6200 ;
  END
END OAI22_X1M_A12TH

MACRO OAI22_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.5550 ;
        RECT 0.8750 0.3200 0.9650 0.5550 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.0500 0.8400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.2500 1.0750 1.3500 ;
        RECT 0.9750 0.9400 1.0750 1.2500 ;
        RECT 0.2000 0.9300 0.3000 1.2500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 1.2500 2.1150 1.3500 ;
        RECT 1.2400 1.0000 1.3400 1.2500 ;
        RECT 2.0150 0.9400 2.1150 1.2500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4700 1.0500 1.8900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7600 2.3500 1.4500 ;
        RECT 0.6100 1.4500 2.3500 1.5500 ;
        RECT 1.3350 0.6600 2.3500 0.7600 ;
        RECT 0.6100 1.5500 0.7100 1.8750 ;
        RECT 1.6500 1.5500 1.7500 1.8750 ;
    END
    ANTENNADIFFAREA 0.426 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.1350 1.6600 1.2250 2.0800 ;
        RECT 2.1750 1.6600 2.2650 2.0800 ;
        RECT 0.0950 1.6400 0.1850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1350 0.4800 2.3250 0.5700 ;
      RECT 0.0900 0.6950 1.2250 0.7850 ;
      RECT 1.1350 0.5700 1.2250 0.6950 ;
      RECT 0.0900 0.4100 0.1800 0.6950 ;
      RECT 0.6150 0.4100 0.7050 0.6950 ;
  END
END OAI22_X1P4M_A12TH

MACRO OAI22_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6400 ;
        RECT 0.8750 0.3200 0.9650 0.6400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7600 2.3500 1.4500 ;
        RECT 0.6100 1.4500 2.3500 1.5500 ;
        RECT 1.3350 0.6600 2.3500 0.7600 ;
        RECT 0.6100 1.5500 0.7100 1.8600 ;
        RECT 1.6500 1.5500 1.7500 1.8600 ;
    END
    ANTENNADIFFAREA 0.6 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4750 1.0500 1.8950 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2350 1.2500 2.1150 1.3500 ;
        RECT 1.2350 0.9650 1.3350 1.2500 ;
        RECT 2.0150 0.9650 2.1150 1.2500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1700 1.2500 1.0750 1.3500 ;
        RECT 0.1700 0.9950 0.2700 1.2500 ;
        RECT 0.9750 0.9650 1.0750 1.2500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.0500 0.8550 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0950 1.7900 0.1850 2.0800 ;
        RECT 1.1350 1.7900 1.2250 2.0800 ;
        RECT 2.1750 1.7900 2.2650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1350 0.4800 2.3250 0.5700 ;
      RECT 0.0900 0.7350 1.2250 0.8250 ;
      RECT 1.1350 0.5700 1.2250 0.7350 ;
      RECT 0.0900 0.4100 0.1800 0.7350 ;
      RECT 0.6150 0.4100 0.7050 0.7350 ;
  END
END OAI22_X2M_A12TH

MACRO OA22_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6800 ;
        RECT 1.3700 0.3200 1.4600 0.8900 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0150 0.1600 1.4000 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9900 0.5600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8300 1.1800 1.1900 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.0800 1.6400 0.1700 2.0800 ;
        RECT 1.1200 1.6000 1.2100 2.0800 ;
        RECT 1.3700 1.5950 1.4600 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0100 0.7700 1.3600 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9700 1.7500 1.4400 ;
        RECT 1.6300 1.4400 1.7500 1.8700 ;
        RECT 1.6300 0.5600 1.7500 0.9700 ;
    END
    ANTENNADIFFAREA 0.1848 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.6000 0.4800 1.2100 0.5700 ;
      RECT 1.1200 0.5700 1.2100 0.7100 ;
      RECT 0.0800 0.8000 0.6900 0.8900 ;
      RECT 0.6000 0.5700 0.6900 0.8000 ;
      RECT 0.0800 0.4800 0.1700 0.8000 ;
      RECT 0.8600 1.3100 1.5450 1.4000 ;
      RECT 1.4550 1.0700 1.5450 1.3100 ;
      RECT 0.5600 1.7900 0.7300 1.9900 ;
      RECT 0.5600 1.7000 0.9500 1.7900 ;
      RECT 0.8600 1.4000 0.9500 1.7000 ;
      RECT 0.8600 0.6900 0.9500 1.3100 ;
  END
END OA22_X0P7M_A12TH

MACRO OA22_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.5950 ;
        RECT 1.3700 0.3200 1.4600 0.6650 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1600 1.3950 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0100 0.5600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0100 1.1600 1.3950 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.3700 1.7700 1.4600 2.0800 ;
        RECT 0.0800 1.7300 0.1700 2.0800 ;
        RECT 1.1200 1.7300 1.2100 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0100 0.7700 1.3600 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9600 1.7500 1.2900 ;
        RECT 1.6300 1.2900 1.7500 1.7200 ;
        RECT 1.6300 0.5500 1.7500 0.9600 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8000 0.6900 0.8900 ;
      RECT 0.6000 0.5700 0.6900 0.8000 ;
      RECT 0.6000 0.4800 1.2100 0.5700 ;
      RECT 1.1200 0.5700 1.2100 0.8900 ;
      RECT 0.0800 0.4600 0.1700 0.8000 ;
      RECT 0.8600 1.5200 1.5300 1.6100 ;
      RECT 1.4400 1.0300 1.5300 1.5200 ;
      RECT 0.5600 1.7700 0.7300 1.9700 ;
      RECT 0.5600 1.6800 0.9500 1.7700 ;
      RECT 0.8600 1.6100 0.9500 1.6800 ;
      RECT 0.8600 0.6900 0.9500 1.5200 ;
  END
END OA22_X1M_A12TH

MACRO OA22_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.4300 0.3200 0.5200 0.6100 ;
        RECT 2.1100 0.3200 2.2000 0.8900 ;
        RECT 2.6300 0.3200 2.7200 0.8900 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3700 1.4500 2.7550 1.5500 ;
        RECT 2.3700 1.5500 2.4600 1.9650 ;
        RECT 2.6650 1.0900 2.7550 1.4500 ;
        RECT 2.3700 1.0000 2.7550 1.0900 ;
        RECT 2.3700 0.5400 2.4600 1.0000 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5200 1.0500 1.8950 1.1950 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3800 1.4500 2.0950 1.5400 ;
        RECT 1.8100 1.5400 2.0950 1.5500 ;
        RECT 1.3800 1.4450 1.4700 1.4500 ;
        RECT 2.0050 1.2950 2.0950 1.4500 ;
        RECT 1.2600 1.3550 1.4700 1.4450 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.0500 0.7900 1.2000 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.4750 0.9700 1.5500 ;
        RECT 0.1550 1.4500 0.9700 1.4750 ;
        RECT 0.1550 1.3850 0.3650 1.4500 ;
        RECT 0.8800 1.0650 0.9700 1.4500 ;
        RECT 0.8800 0.9750 1.1100 1.0650 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.1500 1.8200 1.2400 2.0800 ;
        RECT 2.1100 1.8200 2.2000 2.0800 ;
        RECT 0.1200 1.7500 0.2100 2.0800 ;
        RECT 2.6300 1.7500 2.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8100 0.5550 0.9000 ;
      RECT 0.4650 0.8000 0.5550 0.8100 ;
      RECT 0.4650 0.7100 0.9150 0.8000 ;
      RECT 0.7450 0.5750 0.9150 0.7100 ;
      RECT 0.7450 0.4850 1.7550 0.5750 ;
      RECT 1.1050 0.5750 1.2750 0.7750 ;
      RECT 1.6650 0.5750 1.7550 0.9000 ;
      RECT 0.0800 0.4850 0.1700 0.8100 ;
      RECT 2.1850 1.2500 2.5750 1.3400 ;
      RECT 0.5600 1.6400 2.2750 1.7300 ;
      RECT 2.1850 1.3400 2.2750 1.6400 ;
      RECT 0.5600 1.7300 0.7300 1.9300 ;
      RECT 1.0800 1.2450 1.1700 1.6400 ;
      RECT 1.0800 1.1550 1.3100 1.2450 ;
      RECT 1.2200 0.9550 1.3100 1.1550 ;
      RECT 1.6050 1.7300 1.7750 1.9300 ;
      RECT 1.2200 0.8650 1.5350 0.9550 ;
      RECT 1.3650 0.6650 1.5350 0.8650 ;
  END
END OA22_X1P4M_A12TH

MACRO OA22_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.7100 ;
        RECT 0.8600 0.3200 0.9500 0.7100 ;
        RECT 2.4600 0.3200 2.6300 0.5600 ;
        RECT 3.0200 0.3200 3.1100 0.6650 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1850 1.2500 1.0650 1.3500 ;
        RECT 0.1850 1.0400 0.2850 1.2500 ;
        RECT 0.9650 1.0400 1.0650 1.2500 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 1.0500 0.8350 1.1500 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2650 1.2500 2.1500 1.3500 ;
        RECT 1.2650 1.0400 1.3650 1.2500 ;
        RECT 2.0500 1.0400 2.1500 1.2500 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.5000 1.7700 2.5900 2.0800 ;
        RECT 3.0200 1.7700 3.1100 2.0800 ;
        RECT 0.0800 1.6850 0.1700 2.0800 ;
        RECT 1.1200 1.6850 1.2100 2.0800 ;
        RECT 2.1600 1.6850 2.2500 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4850 1.0500 1.9150 1.1600 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9500 3.1500 1.3000 ;
        RECT 2.7550 1.3000 3.1500 1.4000 ;
        RECT 2.7550 0.8500 3.1500 0.9500 ;
        RECT 2.7550 1.4000 2.8550 1.7300 ;
        RECT 2.7550 0.5400 2.8550 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8300 1.2100 0.9200 ;
      RECT 1.1200 0.5700 1.2100 0.8300 ;
      RECT 1.1200 0.4800 2.3100 0.5700 ;
      RECT 0.0800 0.4600 0.1700 0.8300 ;
      RECT 0.6000 0.4600 0.6900 0.8300 ;
      RECT 2.5000 1.0900 2.9300 1.1800 ;
      RECT 0.6000 1.5000 2.5900 1.5900 ;
      RECT 2.5000 1.1800 2.5900 1.5000 ;
      RECT 2.5000 0.7600 2.5900 1.0900 ;
      RECT 1.3200 0.6700 2.5900 0.7600 ;
      RECT 1.6400 1.5900 1.7300 1.9300 ;
      RECT 0.6000 1.5900 0.6900 1.9300 ;
  END
END OA22_X2M_A12TH

MACRO OA22_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6350 ;
        RECT 0.8600 0.3200 0.9500 0.6350 ;
        RECT 1.1100 0.3200 1.2000 0.6350 ;
        RECT 3.0500 0.3200 3.1400 0.6750 ;
        RECT 3.5700 0.3200 3.6600 0.6750 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7600 1.1200 1.9500 1.3000 ;
        RECT 1.7600 1.3000 2.7400 1.3200 ;
        RECT 1.7600 1.3200 2.5700 1.3900 ;
        RECT 2.4800 1.2300 2.7400 1.3000 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1150 1.0500 3.0200 1.1400 ;
        RECT 2.1150 1.1400 2.3900 1.2000 ;
        RECT 2.9300 1.1400 3.0200 1.2600 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.1000 0.8350 1.2000 ;
        RECT 0.6100 1.0700 0.8350 1.1000 ;
        RECT 0.6100 0.9800 1.5350 1.0700 ;
        RECT 1.4450 1.0700 1.5350 1.2550 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.2900 1.3000 1.3800 ;
        RECT 0.9650 1.1600 1.3000 1.2900 ;
        RECT 0.2350 1.0850 0.3250 1.2900 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3100 1.2500 3.9200 1.3500 ;
        RECT 3.3100 1.3500 3.4000 1.7200 ;
        RECT 3.8300 1.3500 3.9200 1.7200 ;
        RECT 3.8300 0.9800 3.9200 1.2500 ;
        RECT 3.3100 0.8900 3.9200 0.9800 ;
        RECT 3.3100 0.5300 3.4000 0.8900 ;
        RECT 3.8300 0.5300 3.9200 0.8900 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 3.5700 1.7700 3.6600 2.0800 ;
        RECT 0.1050 1.7500 0.1950 2.0800 ;
        RECT 1.0900 1.7500 1.1800 2.0800 ;
        RECT 2.1150 1.7500 2.2050 2.0800 ;
        RECT 3.0500 1.7500 3.1400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7450 1.7200 0.8350 ;
      RECT 1.6300 0.5700 1.7200 0.7450 ;
      RECT 1.3700 0.4100 1.4600 0.7450 ;
      RECT 1.6300 0.4800 2.7600 0.5700 ;
      RECT 2.1500 0.5700 2.2400 0.7800 ;
      RECT 2.6700 0.5700 2.7600 0.7800 ;
      RECT 1.6300 0.4200 1.7200 0.4800 ;
      RECT 2.1500 0.4100 2.2400 0.4800 ;
      RECT 2.6700 0.4100 2.7600 0.4800 ;
      RECT 0.0800 0.4100 0.1700 0.7450 ;
      RECT 0.6000 0.4100 0.6900 0.7450 ;
      RECT 3.1100 1.0700 3.6050 1.1600 ;
      RECT 0.6000 1.5900 0.6900 1.9300 ;
      RECT 1.6000 1.5900 1.6900 1.9300 ;
      RECT 1.8500 0.6650 2.0200 0.8700 ;
      RECT 2.5900 1.5900 2.6800 1.9200 ;
      RECT 2.3700 0.6650 2.5400 0.8700 ;
      RECT 0.6000 1.5000 3.2000 1.5900 ;
      RECT 3.1100 1.1600 3.2000 1.5000 ;
      RECT 3.1100 0.9600 3.2000 1.0700 ;
      RECT 1.8500 0.8700 3.2000 0.9600 ;
  END
END OA22_X3M_A12TH

MACRO OA22_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6800 ;
        RECT 0.8600 0.3200 0.9500 0.6800 ;
        RECT 1.3800 0.3200 1.4700 0.6800 ;
        RECT 1.6300 0.3200 1.7200 0.7100 ;
        RECT 4.1900 0.3200 4.2800 0.6750 ;
        RECT 4.7100 0.3200 4.8000 0.6750 ;
        RECT 5.2300 0.3200 5.3200 0.6750 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.0250 2.0550 1.1150 ;
        RECT 0.2350 1.1150 0.3250 1.2350 ;
        RECT 1.0100 1.1150 1.3800 1.1500 ;
        RECT 1.9650 1.1150 2.0550 1.2350 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3450 1.0600 4.1200 1.1500 ;
        RECT 2.3450 1.1500 2.5300 1.1650 ;
        RECT 3.1600 1.0450 4.1200 1.0600 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.2400 1.8550 1.3500 ;
        RECT 0.4650 1.2050 0.8350 1.2400 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.2750 3.8350 1.3400 ;
        RECT 2.8100 1.3400 3.8350 1.3650 ;
        RECT 2.6400 1.2400 3.0200 1.2750 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4100 1.2500 5.1850 1.3500 ;
        RECT 4.4100 1.3500 4.5800 1.6300 ;
        RECT 4.9700 1.3500 5.0600 1.7250 ;
        RECT 5.0950 0.9800 5.1850 1.2500 ;
        RECT 4.4500 0.8900 5.1850 0.9800 ;
        RECT 4.4500 0.5300 4.5400 0.8900 ;
        RECT 4.9700 0.5300 5.0600 0.8900 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 0.1300 1.7700 0.2200 2.0800 ;
        RECT 1.1300 1.7700 1.2200 2.0800 ;
        RECT 2.1950 1.7700 2.2850 2.0800 ;
        RECT 3.2450 1.7700 3.3350 2.0800 ;
        RECT 4.1900 1.7700 4.2800 2.0800 ;
        RECT 4.7100 1.7700 4.8000 2.0800 ;
        RECT 5.2300 1.7700 5.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8000 1.9800 0.8900 ;
      RECT 1.8900 0.5700 1.9800 0.8000 ;
      RECT 1.8900 0.4800 3.9800 0.5700 ;
      RECT 2.1900 0.5700 2.3600 0.7700 ;
      RECT 2.7100 0.5700 2.8800 0.7700 ;
      RECT 3.2650 0.5700 3.4350 0.7700 ;
      RECT 3.8100 0.5700 3.9800 0.7700 ;
      RECT 0.0800 0.4600 0.1700 0.8000 ;
      RECT 0.6000 0.4600 0.6900 0.8000 ;
      RECT 1.1200 0.4600 1.2100 0.8000 ;
      RECT 4.2300 1.0700 4.9850 1.1600 ;
      RECT 0.6000 1.5900 0.6900 1.9300 ;
      RECT 1.6300 1.5900 1.7200 1.9300 ;
      RECT 2.1450 0.9550 2.2350 1.5000 ;
      RECT 0.6000 1.5000 2.8400 1.5900 ;
      RECT 2.7500 1.5900 2.8400 1.9300 ;
      RECT 2.9700 0.6600 3.1400 0.8650 ;
      RECT 2.4500 0.6600 2.6200 0.8650 ;
      RECT 3.5500 0.6600 3.7200 0.8650 ;
      RECT 3.7050 1.5900 3.7950 1.9300 ;
      RECT 2.1450 0.8650 4.3200 0.9550 ;
      RECT 4.2300 0.9550 4.3200 1.0700 ;
      RECT 4.2300 1.1600 4.3200 1.5000 ;
      RECT 3.7050 1.5000 4.3200 1.5900 ;
  END
END OA22_X4M_A12TH

MACRO OA22_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6500 ;
        RECT 0.6000 0.3200 0.6900 0.6500 ;
        RECT 1.1200 0.3200 1.2100 0.6500 ;
        RECT 1.6400 0.3200 1.7300 0.5800 ;
        RECT 4.7500 0.3200 4.8400 0.6600 ;
        RECT 5.0100 0.3200 5.1000 0.6600 ;
        RECT 5.5300 0.3200 5.6200 0.6600 ;
        RECT 6.0500 0.3200 6.1400 0.6600 ;
        RECT 6.5700 0.3200 6.6600 0.6600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 1.4750 1.3400 ;
        RECT 0.3350 1.3400 1.4750 1.3500 ;
        RECT 0.2500 0.9550 0.3500 1.2500 ;
        RECT 0.3350 1.3500 0.4350 1.6350 ;
        RECT 0.8550 1.3500 0.9550 1.6350 ;
        RECT 1.3750 1.3500 1.4750 1.6350 ;
        RECT 0.2500 0.8650 1.4750 0.9550 ;
        RECT 0.3350 0.8550 1.4750 0.8650 ;
        RECT 0.3350 0.5050 0.4350 0.8550 ;
        RECT 0.8550 0.5050 0.9550 0.8550 ;
        RECT 1.3750 0.5050 1.4750 0.8550 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 0.8500 3.5750 0.9400 ;
        RECT 3.4850 0.9400 3.5750 1.0750 ;
        RECT 1.7950 0.9400 2.8950 0.9500 ;
        RECT 3.4850 1.0750 3.9350 1.1650 ;
        RECT 1.7950 0.9500 1.8850 1.1950 ;
        RECT 2.5250 0.9500 2.8950 1.1550 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1250 1.0250 5.4950 1.1500 ;
        RECT 4.4150 0.9350 6.1950 1.0250 ;
        RECT 6.1050 1.0250 6.1950 1.0600 ;
        RECT 4.4150 1.0250 4.5050 1.2300 ;
        RECT 6.1050 1.0600 6.5350 1.1500 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 1.2550 4.1450 1.3500 ;
        RECT 3.0250 1.1350 3.3950 1.2550 ;
        RECT 2.0100 1.1000 2.4050 1.2550 ;
        RECT 4.0550 1.0750 4.1450 1.2550 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8300 1.2600 6.7650 1.3500 ;
        RECT 4.8300 1.2500 6.0150 1.2600 ;
        RECT 6.6750 1.0350 6.7650 1.2600 ;
        RECT 4.8300 1.2050 4.9200 1.2500 ;
        RECT 5.6450 1.1150 6.0150 1.2500 ;
        RECT 4.6600 1.1150 4.9200 1.2050 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
        RECT 1.1200 1.7700 1.2100 2.0800 ;
        RECT 1.6400 1.7700 1.7300 2.0800 ;
        RECT 2.6700 1.7700 2.7600 2.0800 ;
        RECT 3.7100 1.7700 3.8000 2.0800 ;
        RECT 4.7500 1.7700 4.8400 2.0800 ;
        RECT 5.7900 1.7700 5.8800 2.0800 ;
        RECT 6.8300 1.7700 6.9200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.2300 1.5050 6.4000 1.5950 ;
      RECT 6.3100 1.5950 6.4000 1.9300 ;
      RECT 1.6150 0.7600 1.7050 1.0650 ;
      RECT 0.6350 1.0650 1.7050 1.1550 ;
      RECT 1.6150 1.1550 1.7050 1.5000 ;
      RECT 2.1500 1.5900 2.2400 1.9300 ;
      RECT 1.6150 1.5000 3.2800 1.5900 ;
      RECT 3.1900 1.5900 3.2800 1.9300 ;
      RECT 4.2300 1.5950 4.3200 1.9300 ;
      RECT 4.2350 0.7600 4.3250 1.5050 ;
      RECT 1.6150 0.6700 4.3250 0.7600 ;
      RECT 5.2700 1.5950 5.3600 1.9300 ;
      RECT 4.4900 0.7550 6.9200 0.8450 ;
      RECT 6.8300 0.4150 6.9200 0.7550 ;
      RECT 4.4900 0.5700 4.5800 0.7550 ;
      RECT 2.0900 0.4800 4.5800 0.5700 ;
      RECT 4.4900 0.4750 4.5800 0.4800 ;
      RECT 5.2700 0.4150 5.3600 0.7550 ;
      RECT 5.7900 0.4150 5.8800 0.7550 ;
      RECT 6.3100 0.4150 6.4000 0.7550 ;
  END
END OA22_X6M_A12TH

MACRO OA22_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 9.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6500 ;
        RECT 0.6000 0.3200 0.6900 0.6500 ;
        RECT 1.1200 0.3200 1.2100 0.6500 ;
        RECT 1.6400 0.3200 1.7300 0.6500 ;
        RECT 2.1600 0.3200 2.2500 0.5800 ;
        RECT 6.0800 0.3200 6.2500 0.5800 ;
        RECT 6.3700 0.3200 6.4600 0.5800 ;
        RECT 6.8900 0.3200 6.9800 0.5800 ;
        RECT 7.4100 0.3200 7.5000 0.5800 ;
        RECT 7.9300 0.3200 8.0200 0.5800 ;
        RECT 8.4500 0.3200 8.5400 0.5800 ;
        RECT 8.9700 0.3200 9.0600 0.5800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2350 1.9950 1.3550 ;
        RECT 0.3350 1.3550 1.9950 1.3650 ;
        RECT 0.2500 0.9000 0.3500 1.2350 ;
        RECT 0.3350 1.3650 0.4350 1.7200 ;
        RECT 0.8550 1.3650 0.9550 1.7200 ;
        RECT 1.3750 1.3650 1.4750 1.7200 ;
        RECT 1.8950 1.3650 1.9950 1.7200 ;
        RECT 0.2500 0.7700 1.9950 0.9000 ;
        RECT 0.3350 0.4700 0.4350 0.7700 ;
        RECT 0.8550 0.4700 0.9550 0.7700 ;
        RECT 1.3750 0.4700 1.4750 0.7700 ;
        RECT 1.8950 0.4700 1.9950 0.7700 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2650 0.8500 2.7050 0.9250 ;
        RECT 2.2650 0.9250 5.2950 1.0150 ;
        RECT 2.2650 1.0150 3.2250 1.0300 ;
        RECT 3.9050 1.0150 4.2750 1.0750 ;
        RECT 4.9250 1.0150 5.2950 1.0350 ;
        RECT 2.2650 1.0300 2.3550 1.2150 ;
    END
    ANTENNAGATEAREA 0.5985 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0950 0.8550 6.7900 0.9450 ;
        RECT 6.0950 0.9450 6.1900 0.9650 ;
        RECT 6.4950 0.9450 6.7900 0.9650 ;
        RECT 6.6100 0.8500 6.7900 0.8550 ;
        RECT 5.7850 0.9650 6.1900 1.0550 ;
        RECT 6.4950 0.9650 8.9350 1.0550 ;
        RECT 5.7850 1.0550 5.8750 1.2150 ;
        RECT 6.4950 1.0550 6.8650 1.0650 ;
    END
    ANTENNAGATEAREA 0.5985 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4850 1.2550 2.9050 1.3500 ;
        RECT 2.4850 1.1650 5.5150 1.2550 ;
        RECT 5.4250 1.2550 5.5150 1.3050 ;
        RECT 2.4850 1.1550 2.8550 1.1650 ;
        RECT 3.3950 1.1050 3.7650 1.1650 ;
        RECT 4.4250 1.1050 4.7950 1.1650 ;
        RECT 5.4250 1.0950 5.5150 1.1650 ;
    END
    ANTENNAGATEAREA 0.5985 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4150 1.2550 7.3000 1.3500 ;
        RECT 6.4150 1.2500 9.1650 1.2550 ;
        RECT 6.4150 1.2450 6.5200 1.2500 ;
        RECT 7.0100 1.1550 9.1650 1.2500 ;
        RECT 6.0050 1.1550 6.5200 1.2450 ;
        RECT 9.0750 1.0050 9.1650 1.1550 ;
    END
    ANTENNAGATEAREA 0.5985 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 9.4450 2.7200 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
        RECT 1.1200 1.7700 1.2100 2.0800 ;
        RECT 1.6400 1.7700 1.7300 2.0800 ;
        RECT 2.1600 1.7700 2.2500 2.0800 ;
        RECT 3.0900 1.7500 3.1800 2.0800 ;
        RECT 4.0500 1.7500 4.1400 2.0800 ;
        RECT 5.0600 1.7500 5.1500 2.0800 ;
        RECT 6.1300 1.7500 6.2200 2.0800 ;
        RECT 7.1500 1.7500 7.2400 2.0800 ;
        RECT 8.1900 1.7500 8.2800 2.0800 ;
        RECT 9.2100 1.7500 9.3000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 5.6000 1.5000 8.8000 1.5900 ;
      RECT 8.7100 1.5900 8.8000 1.9300 ;
      RECT 2.0850 1.1350 2.1750 1.5000 ;
      RECT 0.6600 1.0450 2.1750 1.1350 ;
      RECT 2.0850 0.7600 2.1750 1.0450 ;
      RECT 2.6250 1.5900 2.7150 1.9300 ;
      RECT 3.5600 1.5900 3.6500 1.9300 ;
      RECT 2.0850 1.5000 4.6600 1.5900 ;
      RECT 4.5700 1.5900 4.6600 1.9300 ;
      RECT 2.0850 0.6700 5.6950 0.7600 ;
      RECT 5.6050 0.7600 5.6950 1.4650 ;
      RECT 5.6000 1.4650 5.6950 1.5000 ;
      RECT 5.6000 1.5900 5.6900 1.9300 ;
      RECT 6.6300 1.5900 6.7200 1.9300 ;
      RECT 7.6700 1.5900 7.7600 1.9300 ;
      RECT 5.8600 0.6900 9.3200 0.7600 ;
      RECT 7.1500 0.7600 9.3200 0.7800 ;
      RECT 9.2300 0.4100 9.3200 0.6900 ;
      RECT 5.8600 0.7600 5.9500 0.7800 ;
      RECT 5.8600 0.5700 5.9500 0.6700 ;
      RECT 2.4300 0.4800 5.9500 0.5700 ;
      RECT 5.8600 0.4100 5.9500 0.4800 ;
      RECT 6.6300 0.4800 6.7200 0.6700 ;
      RECT 5.8600 0.6700 7.2400 0.6900 ;
      RECT 7.1500 0.4100 7.2400 0.6700 ;
      RECT 7.6700 0.4100 7.7600 0.6900 ;
      RECT 8.1900 0.4100 8.2800 0.6900 ;
      RECT 8.7100 0.4100 8.8000 0.6900 ;
  END
END OA22_X8M_A12TH

MACRO OAI211_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.5300 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8200 0.5600 1.2100 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 0.8100 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7950 1.1600 1.1900 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6450 1.3500 1.3000 ;
        RECT 0.6300 1.3000 1.3500 1.4000 ;
        RECT 1.0950 0.5550 1.3500 0.6450 ;
        RECT 0.6300 1.4000 0.7300 1.7200 ;
        RECT 1.1600 1.4000 1.2500 1.7200 ;
    END
    ANTENNADIFFAREA 0.198925 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9000 1.5100 0.9900 2.0800 ;
        RECT 0.1050 1.3400 0.1950 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 0.8200 0.9500 1.2100 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.1050 0.6300 0.7250 0.7200 ;
      RECT 0.6350 0.4950 0.7250 0.6300 ;
      RECT 0.1050 0.4950 0.1950 0.6300 ;
  END
END OAI211_X0P5M_A12TH

MACRO OAI211_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4000 0.3200 0.4900 0.6850 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9950 0.3500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8300 1.0200 0.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9400 1.1500 1.3700 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8300 1.3500 1.5000 ;
        RECT 0.6700 1.5000 1.3500 1.5900 ;
        RECT 1.2050 0.4400 1.3500 0.8300 ;
        RECT 0.6700 1.5900 0.7600 1.8500 ;
        RECT 1.2150 1.5900 1.3050 1.8500 ;
    END
    ANTENNADIFFAREA 0.253525 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9550 1.7500 1.0450 2.0800 ;
        RECT 0.1350 1.5300 0.2250 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0000 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.1350 0.8000 0.7600 0.8900 ;
      RECT 0.6700 0.4450 0.7600 0.8000 ;
      RECT 0.1350 0.4450 0.2250 0.8000 ;
  END
END OAI211_X0P7M_A12TH

MACRO OAI211_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6300 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1600 1.4400 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0100 0.9500 1.3950 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.5600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.8650 1.8600 1.0350 2.0800 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9000 1.3500 1.6500 ;
        RECT 0.6150 1.6500 1.3500 1.7500 ;
        RECT 1.1700 0.4900 1.3500 0.9000 ;
        RECT 0.6150 1.7500 0.7050 1.9600 ;
        RECT 1.1700 1.7500 1.2600 1.9600 ;
    END
    ANTENNADIFFAREA 0.3574 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0450 1.1300 1.1550 1.5400 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END C0
  OBS
    LAYER M1 ;
      RECT 0.0950 0.8100 0.7050 0.9000 ;
      RECT 0.6150 0.4700 0.7050 0.8100 ;
      RECT 0.0950 0.4700 0.1850 0.8100 ;
  END
END OAI211_X1M_A12TH

MACRO OAI211_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7600 ;
        RECT 0.8750 0.3200 0.9650 0.7600 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.2500 1.0800 1.3500 ;
        RECT 0.1950 1.1400 0.2950 1.2500 ;
        RECT 0.9800 1.1400 1.0800 1.2500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2550 1.2500 2.1400 1.3500 ;
        RECT 1.2550 1.1400 1.3550 1.2500 ;
        RECT 2.0400 1.1400 2.1400 1.2500 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 1.0500 1.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END C0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.6400 1.6700 1.8100 2.0800 ;
        RECT 2.1750 1.6700 2.3450 2.0800 ;
        RECT 0.0950 1.6550 0.1850 2.0800 ;
        RECT 1.0850 1.6550 1.1750 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.4500 ;
        RECT 0.6100 1.4500 2.3500 1.5500 ;
        RECT 1.6800 0.8500 2.3500 0.9500 ;
        RECT 0.6100 1.5500 0.7100 1.9050 ;
        RECT 1.4200 1.5500 1.5100 1.6900 ;
        RECT 1.9400 1.5500 2.0300 1.6900 ;
        RECT 1.6800 0.7150 1.7700 0.8500 ;
    END
    ANTENNADIFFAREA 0.3638 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.1350 0.4800 2.3550 0.5700 ;
      RECT 0.0950 0.8550 1.2250 0.9450 ;
      RECT 1.1350 0.5700 1.2250 0.8550 ;
      RECT 0.0950 0.4900 0.1850 0.8550 ;
      RECT 0.6150 0.4950 0.7050 0.8550 ;
  END
END OAI211_X1P4M_A12TH

MACRO OAI211_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6300 ;
        RECT 0.8750 0.3200 0.9650 0.6300 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.2500 1.1250 1.3500 ;
        RECT 0.2450 1.0500 0.3450 1.2500 ;
        RECT 1.0250 1.0500 1.1250 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5100 1.2500 1.9300 1.3500 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3000 1.0500 2.1500 1.1500 ;
        RECT 1.3000 1.1500 1.4000 1.2800 ;
        RECT 2.0500 1.1500 2.1500 1.2700 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.0500 0.9000 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.4500 ;
        RECT 0.6100 1.4500 2.3500 1.5500 ;
        RECT 1.6700 0.8500 2.3500 0.9500 ;
        RECT 0.6100 1.5500 0.7100 1.8800 ;
        RECT 1.4050 1.5500 1.5050 1.9600 ;
        RECT 1.9250 1.5500 2.0250 1.9600 ;
        RECT 1.6700 0.7400 1.7600 0.8500 ;
    END
    ANTENNADIFFAREA 0.515 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 1.6700 1.7700 1.7600 2.0800 ;
        RECT 2.2100 1.7700 2.3000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1350 0.4800 2.3250 0.5700 ;
      RECT 0.0950 0.8100 1.2250 0.9000 ;
      RECT 1.1350 0.5700 1.2250 0.8100 ;
      RECT 0.0950 0.4700 0.1850 0.8100 ;
      RECT 0.6150 0.4700 0.7050 0.8100 ;
  END
END OAI211_X2M_A12TH

MACRO OAI211_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6300 ;
        RECT 0.8750 0.3200 0.9650 0.6300 ;
        RECT 1.3950 0.3200 1.4850 0.6300 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2700 1.0500 0.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0700 1.0500 1.6050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0500 2.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.0500 3.1250 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.5700 3.3500 1.2500 ;
        RECT 1.1350 1.2500 3.3500 1.3500 ;
        RECT 2.6350 0.4800 3.3500 0.5700 ;
        RECT 1.1350 1.3500 1.2250 1.7300 ;
        RECT 1.6550 1.3500 1.7450 1.7700 ;
        RECT 2.1750 1.3500 2.2650 1.7700 ;
        RECT 2.6950 1.3500 2.7850 1.7700 ;
        RECT 3.2150 1.3500 3.3050 1.7700 ;
    END
    ANTENNADIFFAREA 0.85665 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 0.6150 1.7700 0.7050 2.0800 ;
        RECT 1.8750 1.4700 2.0450 2.0800 ;
        RECT 2.3950 1.4700 2.5650 2.0800 ;
        RECT 2.9150 1.4700 3.0850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 0.8300 1.7450 0.9200 ;
      RECT 1.6550 0.5700 1.7450 0.8300 ;
      RECT 1.6550 0.4800 2.3250 0.5700 ;
      RECT 0.0950 0.4900 0.1850 0.8300 ;
      RECT 0.6150 0.4900 0.7050 0.8300 ;
      RECT 1.1350 0.4900 1.2250 0.8300 ;
      RECT 1.8550 0.7700 3.1050 0.8600 ;
      RECT 2.4350 0.4300 2.5250 0.7700 ;
      RECT 0.8750 1.8300 1.4850 1.9200 ;
      RECT 1.3950 1.4900 1.4850 1.8300 ;
      RECT 0.3550 1.4800 0.9650 1.5700 ;
      RECT 0.8750 1.5700 0.9650 1.8300 ;
      RECT 0.3550 1.5700 0.4450 1.9100 ;
  END
END OAI211_X3M_A12TH

MACRO OAI211_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6300 ;
        RECT 0.8750 0.3200 0.9650 0.6300 ;
        RECT 1.3950 0.3200 1.4850 0.6300 ;
        RECT 1.9150 0.3200 2.0050 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 2.7800 1.7850 2.8700 2.0800 ;
        RECT 3.3000 1.7850 3.3900 2.0800 ;
        RECT 3.8200 1.7850 3.9100 2.0800 ;
        RECT 4.3400 1.7850 4.4300 2.0800 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 2.2050 1.7700 2.2950 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9500 4.5500 1.4500 ;
        RECT 0.6150 1.4500 4.5500 1.5500 ;
        RECT 2.7800 0.8500 4.5500 0.9500 ;
        RECT 0.6150 1.5500 0.7050 1.8800 ;
        RECT 1.6550 1.5500 1.7450 1.8800 ;
        RECT 2.5200 1.5500 2.6100 1.9600 ;
        RECT 3.0400 1.5500 3.1300 1.9600 ;
        RECT 3.5600 1.5500 3.6500 1.9600 ;
        RECT 4.0800 1.5500 4.1700 1.9600 ;
        RECT 2.7800 0.7400 2.8700 0.8500 ;
        RECT 3.8200 0.7400 3.9100 0.8500 ;
    END
    ANTENNADIFFAREA 1.012 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6450 1.2500 4.0950 1.3500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END C0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0550 2.1500 1.2600 ;
        RECT 0.2450 0.9550 2.1500 1.0550 ;
        RECT 0.2450 1.0550 0.3450 1.2600 ;
        RECT 1.0100 1.0550 1.4100 1.1500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.2550 1.6200 1.3500 ;
        RECT 0.4800 1.2500 1.9300 1.2550 ;
        RECT 0.4800 1.1550 0.8900 1.2500 ;
        RECT 1.5200 1.1550 1.9300 1.2500 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4100 1.0500 4.3300 1.1500 ;
        RECT 2.4100 1.1500 2.5100 1.3250 ;
        RECT 4.2300 1.1500 4.3300 1.2800 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 2.2300 0.4800 4.4900 0.5700 ;
      RECT 0.0950 0.7600 2.3200 0.8500 ;
      RECT 2.2300 0.5700 2.3200 0.7600 ;
      RECT 0.0950 0.4300 0.1850 0.7600 ;
      RECT 0.6150 0.4300 0.7050 0.7600 ;
      RECT 1.1350 0.4300 1.2250 0.7600 ;
      RECT 1.6550 0.4300 1.7450 0.7600 ;
  END
END OAI211_X4M_A12TH

MACRO OAI21B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.5600 ;
        RECT 1.2200 0.3200 1.3200 0.9900 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.5050 1.1900 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1950 0.1600 1.5900 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9850 1.2500 1.2550 1.3500 ;
        RECT 1.1450 1.1000 1.2550 1.2500 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END B0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9000 1.7250 1.0700 2.0800 ;
        RECT 0.0750 1.7200 0.1750 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7850 0.4500 1.0100 0.5750 ;
        RECT 0.7850 0.5750 0.8750 0.8500 ;
        RECT 0.5950 0.8500 0.8750 0.9500 ;
        RECT 0.5950 0.9500 0.6950 1.9900 ;
    END
    ANTENNADIFFAREA 0.1547 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0750 0.6500 0.6900 0.7400 ;
      RECT 0.5950 0.5250 0.6900 0.6500 ;
      RECT 0.0750 0.5000 0.1750 0.6500 ;
      RECT 1.2250 1.6250 1.3150 1.8450 ;
      RECT 0.7850 1.5350 1.3150 1.6250 ;
      RECT 0.7850 1.0400 1.0550 1.1300 ;
      RECT 0.9650 0.8100 1.0550 1.0400 ;
      RECT 0.7850 1.1300 0.8750 1.5350 ;
  END
END OAI21B_X0P5M_A12TH

MACRO OAI21B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3700 0.3200 0.4700 0.7100 ;
        RECT 1.4300 0.3200 1.5200 0.9000 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0400 0.5500 1.4250 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6900 1.2900 0.9500 1.3900 ;
        RECT 0.6900 1.3900 0.7900 1.5100 ;
        RECT 0.8500 0.9250 0.9500 1.2900 ;
        RECT 0.6500 1.5100 0.7900 1.7200 ;
        RECT 0.8500 0.5150 1.0000 0.9250 ;
    END
    ANTENNADIFFAREA 0.179075 ;
  END Y

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.2800 1.5500 1.5950 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END B0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.4300 1.7150 1.5200 2.0800 ;
        RECT 0.1100 1.6600 0.2000 2.0800 ;
        RECT 0.9100 1.5700 1.0000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1150 0.8300 0.7250 0.9200 ;
      RECT 0.6350 0.5100 0.7250 0.8300 ;
      RECT 0.1150 0.5100 0.2050 0.8300 ;
      RECT 1.1700 1.2750 1.2600 1.9250 ;
      RECT 1.0700 1.0650 1.2600 1.2750 ;
      RECT 1.1700 0.6900 1.2600 1.0650 ;
  END
END OAI21B_X0P7M_A12TH

MACRO OAI21B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6500 ;
        RECT 1.4300 0.3200 1.5200 0.8800 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9950 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.0500 0.7100 1.1500 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8500 0.9500 1.3000 ;
        RECT 0.6100 1.3000 0.9500 1.4000 ;
        RECT 0.8500 0.4400 1.0000 0.8500 ;
        RECT 0.6100 1.4000 0.7100 1.7300 ;
    END
    ANTENNADIFFAREA 0.26425 ;
  END Y

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.2900 1.5500 1.5900 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END B0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.0950 1.7350 0.1850 2.0800 ;
        RECT 1.4300 1.7100 1.5200 2.0800 ;
        RECT 0.8900 1.5550 0.9800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 0.7700 0.7050 0.8600 ;
      RECT 0.6150 0.4400 0.7050 0.7700 ;
      RECT 0.0950 0.4400 0.1850 0.7700 ;
      RECT 1.1700 1.1800 1.2600 1.9200 ;
      RECT 1.0700 0.9700 1.2600 1.1800 ;
      RECT 1.1700 0.6700 1.2600 0.9700 ;
  END
END OAI21B_X1M_A12TH

MACRO OAI21B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6500 ;
        RECT 0.8600 0.3200 0.9500 0.6500 ;
        RECT 2.2300 0.3200 2.3200 0.7000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.6950 1.5500 1.5200 ;
        RECT 0.6000 1.5200 1.5500 1.6100 ;
        RECT 0.6000 1.6100 0.6900 1.9500 ;
        RECT 1.4500 1.6100 1.5500 1.8050 ;
    END
    ANTENNADIFFAREA 0.28 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0100 1.1500 1.3000 ;
        RECT 0.1850 1.3000 1.1500 1.4000 ;
        RECT 0.1850 1.0100 0.2850 1.3000 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 1.0500 0.8450 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 1.0800 2.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END B0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.1200 1.7100 1.2100 2.0800 ;
        RECT 0.0800 1.6100 0.1700 2.0800 ;
        RECT 1.7150 1.5500 1.8050 2.0800 ;
        RECT 2.2300 1.5100 2.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1600 0.4800 1.8050 0.5700 ;
      RECT 1.7150 0.5700 1.8050 0.8900 ;
      RECT 0.0800 0.8000 1.2500 0.8900 ;
      RECT 1.1600 0.5700 1.2500 0.8000 ;
      RECT 0.0800 0.4500 0.1700 0.8000 ;
      RECT 0.6000 0.4800 0.6900 0.8000 ;
      RECT 1.9700 1.1200 2.0600 1.6650 ;
      RECT 1.6700 1.0300 2.0600 1.1200 ;
      RECT 1.9700 0.4900 2.0600 1.0300 ;
  END
END OAI21B_X1P4M_A12TH

MACRO OAI21B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6450 ;
        RECT 0.8750 0.3200 0.9650 0.6450 ;
        RECT 2.2250 0.3200 2.3150 0.7000 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1850 1.2500 1.2000 1.3500 ;
        RECT 0.1850 0.9750 0.3000 1.2500 ;
        RECT 1.1000 0.9750 1.2000 1.2500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.6900 1.5500 1.4500 ;
        RECT 0.6150 1.4500 1.5500 1.5500 ;
        RECT 0.6150 1.5500 0.7050 1.8800 ;
    END
    ANTENNADIFFAREA 0.40865 ;
  END Y

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 0.9950 2.3500 1.2950 ;
    END
    ANTENNAGATEAREA 0.0375 ;
  END B0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 1.1350 1.7700 1.2250 2.0800 ;
        RECT 2.2250 1.5000 2.3150 2.0800 ;
        RECT 1.7150 1.3350 1.8050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1400 0.4800 1.8050 0.5700 ;
      RECT 1.7150 0.5700 1.8050 0.8900 ;
      RECT 0.0800 0.7650 1.2300 0.8550 ;
      RECT 1.1400 0.5700 1.2300 0.7650 ;
      RECT 0.0800 0.4400 0.1700 0.7650 ;
      RECT 0.6000 0.4450 0.6900 0.7650 ;
      RECT 1.9650 1.1150 2.0550 1.8900 ;
      RECT 1.6700 1.0250 2.0550 1.1150 ;
      RECT 1.9650 0.5600 2.0550 1.0250 ;
  END
END OAI21B_X2M_A12TH

MACRO OAI21B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7100 ;
        RECT 0.8750 0.3200 0.9650 0.7100 ;
        RECT 1.3950 0.3200 1.4850 0.7100 ;
        RECT 2.9700 0.3200 3.0600 0.7000 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0500 0.7050 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0800 1.0500 1.5900 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.3450 1.7500 1.7500 ;
        RECT 1.1350 1.2550 2.2900 1.3450 ;
        RECT 1.1350 1.3450 1.2250 1.7000 ;
        RECT 2.1900 1.3450 2.2900 1.7200 ;
        RECT 1.9300 0.7800 2.0200 1.2550 ;
        RECT 1.9300 0.6900 2.5400 0.7800 ;
        RECT 2.4500 0.7800 2.5400 0.9200 ;
        RECT 2.4500 0.5100 2.5400 0.6900 ;
    END
    ANTENNADIFFAREA 0.64155 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0950 1.7700 0.1850 2.0800 ;
        RECT 0.6150 1.7700 0.7050 2.0800 ;
        RECT 2.9700 1.4800 3.0600 2.0800 ;
        RECT 1.8900 1.4600 2.0600 2.0800 ;
        RECT 2.4500 1.3550 2.5400 2.0800 ;
    END
  END VDD

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0300 1.0050 3.1500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0549 ;
  END B0N
  OBS
    LAYER M1 ;
      RECT 2.7100 1.1400 2.8000 1.8100 ;
      RECT 2.1100 1.0500 2.8000 1.1400 ;
      RECT 2.7100 0.5300 2.8000 1.0500 ;
      RECT 0.8750 1.8300 1.4850 1.9200 ;
      RECT 1.3950 1.5100 1.4850 1.8300 ;
      RECT 0.3550 1.5000 0.9650 1.5900 ;
      RECT 0.8750 1.5900 0.9650 1.8300 ;
      RECT 0.3550 1.5900 0.4450 1.9450 ;
      RECT 1.6550 0.4800 2.3400 0.5700 ;
      RECT 0.0950 0.8300 1.7450 0.9200 ;
      RECT 1.6550 0.5700 1.7450 0.8300 ;
      RECT 0.0950 0.4900 0.1850 0.8300 ;
      RECT 0.6150 0.4900 0.7050 0.8300 ;
      RECT 1.1350 0.4900 1.2250 0.8300 ;
  END
END OAI21B_X3M_A12TH

MACRO OAI21B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7100 ;
        RECT 0.8750 0.3200 0.9650 0.7100 ;
        RECT 1.3950 0.3200 1.4850 0.7100 ;
        RECT 1.9150 0.3200 2.0050 0.7100 ;
        RECT 3.7800 0.3200 3.8700 0.8250 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0400 0.9000 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 1.0400 2.0600 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3950 1.2500 3.0500 1.3500 ;
        RECT 1.3950 1.3500 1.4850 1.7000 ;
        RECT 1.9150 1.3500 2.0050 1.7000 ;
        RECT 2.4250 1.3500 2.5250 1.9150 ;
        RECT 2.9500 1.3500 3.0500 1.7200 ;
        RECT 2.4250 0.7900 2.5250 1.2500 ;
        RECT 2.4250 0.6900 3.1150 0.7900 ;
    END
    ANTENNADIFFAREA 0.8286 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 3.7800 1.5800 3.8700 2.0800 ;
        RECT 2.6950 1.4950 2.7850 2.0800 ;
        RECT 3.2200 1.4950 3.3100 2.0800 ;
    END
  END VDD

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.9650 3.7500 1.3850 ;
    END
    ANTENNAGATEAREA 0.0723 ;
  END B0N
  OBS
    LAYER M1 ;
      RECT 1.1350 1.8300 2.2650 1.9200 ;
      RECT 2.1750 1.4900 2.2650 1.8300 ;
      RECT 0.0950 1.5000 1.2250 1.5900 ;
      RECT 1.1350 1.5900 1.2250 1.8300 ;
      RECT 1.6550 1.4900 1.7450 1.8300 ;
      RECT 0.0950 1.5900 0.1850 1.9300 ;
      RECT 0.6150 1.5900 0.7050 1.9300 ;
      RECT 2.1750 0.4800 3.3050 0.5700 ;
      RECT 3.2150 0.5700 3.3050 0.8900 ;
      RECT 0.0950 0.8300 2.2650 0.9200 ;
      RECT 2.1750 0.5700 2.2650 0.8300 ;
      RECT 0.0950 0.4600 0.1850 0.8300 ;
      RECT 0.6150 0.4600 0.7050 0.8300 ;
      RECT 1.1350 0.4600 1.2250 0.8300 ;
      RECT 1.6550 0.4600 1.7450 0.8300 ;
      RECT 3.4600 1.1450 3.5600 1.7650 ;
      RECT 2.6450 1.0550 3.5600 1.1450 ;
      RECT 3.4600 0.4950 3.5600 1.0550 ;
  END
END OAI21B_X4M_A12TH

MACRO OAI21B_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.3700 0.3200 0.4700 0.5450 ;
        RECT 0.8900 0.3200 0.9900 0.5450 ;
        RECT 1.4100 0.3200 1.5100 0.5450 ;
        RECT 1.9300 0.3200 2.0300 0.5450 ;
        RECT 2.4500 0.3200 2.5500 0.5700 ;
        RECT 2.6600 0.3200 2.8350 0.5750 ;
        RECT 4.6650 0.3200 4.7650 0.7800 ;
        RECT 5.1850 0.3200 5.2850 0.8000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 0.1100 1.7700 0.2100 2.0800 ;
        RECT 1.1500 1.7700 1.2500 2.0800 ;
        RECT 2.1900 1.7700 2.2900 2.0800 ;
        RECT 3.1900 1.6450 3.2900 2.0800 ;
        RECT 3.7100 1.6450 3.8100 2.0800 ;
        RECT 4.2300 1.5750 4.3300 2.0800 ;
        RECT 4.6650 1.4400 4.7650 2.0800 ;
        RECT 5.1850 1.4000 5.2850 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0050 1.0500 1.4000 1.1500 ;
        RECT 1.0050 0.9500 1.1050 1.0500 ;
        RECT 1.3000 0.9500 1.4000 1.0500 ;
        RECT 0.2850 0.8500 1.1050 0.9500 ;
        RECT 1.3000 0.8500 2.1500 0.9500 ;
        RECT 0.2850 0.9500 0.3850 1.2100 ;
        RECT 2.0500 0.9500 2.1500 1.0500 ;
        RECT 2.0500 1.0500 2.4300 1.1500 ;
        RECT 2.3300 0.9500 2.4300 1.0500 ;
        RECT 2.3300 0.8500 3.1350 0.9500 ;
        RECT 3.0350 0.9500 3.1350 1.2050 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7950 1.0500 5.2150 1.1500 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END B0N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8300 1.2500 2.6300 1.3500 ;
        RECT 1.8300 1.1650 1.9300 1.2500 ;
        RECT 2.5300 1.1600 2.6300 1.2500 ;
        RECT 1.5200 1.0650 1.9300 1.1650 ;
        RECT 2.5300 1.0600 2.9400 1.1600 ;
        RECT 1.5200 1.1650 1.6200 1.2500 ;
        RECT 0.7700 1.2500 1.6200 1.3500 ;
        RECT 0.7700 1.1700 0.8700 1.2500 ;
        RECT 0.5000 1.0700 0.8700 1.1700 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 1.4500 4.0700 1.5500 ;
        RECT 0.6300 1.5500 0.7300 1.8800 ;
        RECT 1.6700 1.5500 1.7700 1.8250 ;
        RECT 2.6900 1.5500 2.7900 1.8250 ;
        RECT 3.4500 1.5500 3.5500 1.8050 ;
        RECT 3.9700 1.5500 4.0700 1.8800 ;
        RECT 3.3350 1.0000 3.4350 1.4500 ;
        RECT 3.3350 0.9000 4.5050 1.0000 ;
        RECT 3.3350 0.6600 3.5050 0.9000 ;
        RECT 3.8550 0.6600 4.0250 0.9000 ;
        RECT 4.4050 0.5450 4.5050 0.9000 ;
    END
    ANTENNADIFFAREA 1.2296 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 3.0450 0.4800 4.2850 0.5700 ;
      RECT 4.1550 0.5700 4.2850 0.8100 ;
      RECT 0.0750 0.6700 3.1750 0.7600 ;
      RECT 3.0450 0.5700 3.1750 0.6700 ;
      RECT 3.0450 0.4200 3.1750 0.4800 ;
      RECT 3.6350 0.5700 3.7250 0.8100 ;
      RECT 0.0750 0.4200 0.2050 0.6700 ;
      RECT 0.6350 0.4200 0.7250 0.6700 ;
      RECT 1.1550 0.4200 1.2450 0.6700 ;
      RECT 1.6750 0.4200 1.7650 0.6700 ;
      RECT 2.1950 0.4200 2.2850 0.6700 ;
      RECT 4.9300 1.3300 5.0200 1.7500 ;
      RECT 4.5950 1.2400 5.0200 1.3300 ;
      RECT 4.5950 0.8700 5.0200 0.9600 ;
      RECT 4.9300 0.4750 5.0200 0.8700 ;
      RECT 4.5950 1.1800 4.6850 1.2400 ;
      RECT 3.5550 1.0900 4.6850 1.1800 ;
      RECT 4.5950 0.9600 4.6850 1.0900 ;
  END
END OAI21B_X6M_A12TH

MACRO OAI21B_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.8200 ;
        RECT 0.6050 0.3200 0.7050 0.7500 ;
        RECT 3.3750 0.3200 3.4750 0.5700 ;
        RECT 3.8950 0.3200 3.9950 0.5700 ;
        RECT 4.4150 0.3200 4.5150 0.5700 ;
        RECT 4.9350 0.3200 5.0350 0.5700 ;
        RECT 5.4550 0.3200 5.5550 0.5700 ;
        RECT 5.9750 0.3200 6.0750 0.5700 ;
        RECT 6.4950 0.3200 6.5950 0.5700 ;
    END
  END VSS

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.0500 0.5750 1.1600 ;
    END
    ANTENNAGATEAREA 0.1446 ;
  END B0N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3550 0.8500 4.1200 0.9500 ;
        RECT 3.3550 0.9500 3.4550 1.0600 ;
        RECT 4.0200 0.9500 4.1200 0.9600 ;
        RECT 3.0650 1.0600 3.4550 1.1600 ;
        RECT 4.0200 0.9600 4.4100 1.0600 ;
        RECT 4.3100 0.9500 4.4100 0.9600 ;
        RECT 4.3100 0.8500 5.1450 0.9500 ;
        RECT 5.0450 0.9500 5.1450 0.9600 ;
        RECT 5.0450 0.9600 5.4550 1.0600 ;
        RECT 5.3550 0.9500 5.4550 0.9600 ;
        RECT 5.3550 0.9450 6.4650 0.9500 ;
        RECT 6.0450 0.9500 6.4650 1.0450 ;
        RECT 5.3550 0.8500 6.1450 0.9450 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8400 1.2500 4.6250 1.3500 ;
        RECT 3.8400 1.2050 3.9400 1.2500 ;
        RECT 4.5250 1.2050 4.6250 1.2500 ;
        RECT 3.5450 1.1050 3.9400 1.2050 ;
        RECT 4.5250 1.1050 4.9350 1.2050 ;
        RECT 3.5450 1.2050 3.6450 1.2500 ;
        RECT 4.8350 1.2050 4.9350 1.2500 ;
        RECT 2.8300 1.2500 3.6450 1.3500 ;
        RECT 4.8350 1.2500 5.6650 1.3500 ;
        RECT 2.8300 1.0700 2.9300 1.2500 ;
        RECT 5.5650 1.2250 5.6650 1.2500 ;
        RECT 5.5650 1.1250 5.9750 1.2250 ;
        RECT 5.8750 1.2250 5.9750 1.2500 ;
        RECT 5.8750 1.2500 6.6950 1.3500 ;
        RECT 6.5950 0.9800 6.6950 1.2500 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1150 1.4500 6.3250 1.5500 ;
        RECT 1.1150 1.5500 1.2150 1.8600 ;
        RECT 1.6350 1.5500 1.7350 1.8200 ;
        RECT 2.1550 1.5500 2.2550 1.8200 ;
        RECT 3.1950 1.5500 3.2950 1.8200 ;
        RECT 4.1550 1.5500 4.2550 1.8200 ;
        RECT 5.1950 1.5500 5.2950 1.8200 ;
        RECT 6.2250 1.5500 6.3250 1.8800 ;
        RECT 2.2500 0.9650 2.3500 1.4500 ;
        RECT 0.8550 0.8650 2.5150 0.9650 ;
        RECT 1.3750 0.6750 1.4750 0.8650 ;
        RECT 1.8950 0.6750 1.9950 0.8650 ;
        RECT 2.4150 0.6750 2.5150 0.8650 ;
        RECT 0.8550 0.4450 0.9550 0.8650 ;
    END
    ANTENNADIFFAREA 1.7122 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 3.6900 1.7700 3.7900 2.0800 ;
        RECT 4.6750 1.7700 4.7750 2.0800 ;
        RECT 5.7150 1.7700 5.8150 2.0800 ;
        RECT 6.7050 1.7700 6.8050 2.0800 ;
        RECT 1.3750 1.6600 1.4750 2.0800 ;
        RECT 1.8950 1.6500 1.9950 2.0800 ;
        RECT 2.5450 1.6500 2.6450 2.0800 ;
        RECT 0.0850 1.5350 0.1850 2.0800 ;
        RECT 0.6050 1.5350 0.7050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6650 1.0600 2.1250 1.1500 ;
      RECT 0.3500 1.2650 0.7550 1.3550 ;
      RECT 0.6650 1.1500 0.7550 1.2650 ;
      RECT 0.6650 0.9450 0.7550 1.0600 ;
      RECT 0.3500 0.8550 0.7550 0.9450 ;
      RECT 0.3500 1.3550 0.4400 1.7200 ;
      RECT 0.3500 0.4900 0.4400 0.8550 ;
      RECT 2.6800 0.6700 6.8500 0.7600 ;
      RECT 6.7600 0.7600 6.8500 0.8750 ;
      RECT 6.7600 0.4450 6.8500 0.6700 ;
      RECT 2.6800 0.7600 2.7700 0.8500 ;
      RECT 2.6800 0.5700 2.7700 0.6700 ;
      RECT 3.1200 0.4300 3.2100 0.6700 ;
      RECT 1.0800 0.4800 2.7700 0.5700 ;
      RECT 1.0800 0.5700 1.2500 0.7700 ;
      RECT 1.6000 0.5700 1.7700 0.7700 ;
      RECT 2.1200 0.5700 2.2900 0.7700 ;
      RECT 3.6400 0.4300 3.7300 0.6700 ;
      RECT 4.1600 0.4300 4.2500 0.6700 ;
      RECT 4.6800 0.4300 4.7700 0.6700 ;
      RECT 5.2000 0.4300 5.2900 0.6700 ;
      RECT 5.7200 0.4100 5.8100 0.6700 ;
      RECT 6.2400 0.4300 6.3300 0.6700 ;
  END
END OAI21B_X8M_A12TH

MACRO OAI21_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.6950 0.3200 0.7950 0.7400 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9550 0.3500 1.3750 ;
    END
    ANTENNAGATEAREA 0.0321 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.2100 0.7500 1.5650 ;
        RECT 0.5350 1.1100 0.7500 1.2100 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0350 0.9500 1.5050 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7650 0.1500 1.6500 ;
        RECT 0.0500 1.6500 0.5700 1.7500 ;
        RECT 0.0500 0.6650 0.2550 0.7650 ;
        RECT 0.4000 1.7500 0.5700 1.9600 ;
    END
    ANTENNADIFFAREA 0.156725 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.1000 1.8550 0.2000 2.0800 ;
        RECT 0.9550 1.7000 1.0550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4400 0.8300 1.0500 0.9200 ;
      RECT 0.9600 0.6600 1.0500 0.8300 ;
      RECT 0.4400 0.6600 0.5300 0.8300 ;
  END
END OAI21_X0P5M_A12TH

MACRO OAI21_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4100 0.3200 0.5000 0.7250 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0100 0.3550 1.3950 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0100 0.5750 1.3950 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9200 1.1500 1.6500 ;
        RECT 0.6650 1.6500 1.1500 1.7500 ;
        RECT 0.9550 0.8200 1.1500 0.9200 ;
        RECT 0.6650 1.7500 0.7650 1.9650 ;
        RECT 0.9550 0.4900 1.0450 0.8200 ;
    END
    ANTENNADIFFAREA 0.193775 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.0300 0.9500 1.4400 ;
    END
    ANTENNAGATEAREA 0.0453 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9450 1.8800 1.0350 2.0800 ;
        RECT 0.1450 1.6600 0.2350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1500 0.8300 0.7700 0.9200 ;
      RECT 0.6800 0.4900 0.7700 0.8300 ;
      RECT 0.1500 0.4900 0.2400 0.8300 ;
  END
END OAI21_X0P7M_A12TH

MACRO NOR3_X1P4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5600 ;
        RECT 0.5600 0.3200 0.7300 0.5200 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3250 1.4550 1.3950 1.5500 ;
        RECT 0.2350 1.4500 1.5150 1.4550 ;
        RECT 0.2350 1.3650 0.4350 1.4500 ;
        RECT 1.3050 1.3650 1.5150 1.4500 ;
        RECT 0.2350 1.2850 0.3250 1.3650 ;
        RECT 1.4250 1.2850 1.5150 1.3650 ;
    END
    ANTENNAGATEAREA 0.1146 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.8500 0.9900 0.9500 ;
        RECT 0.8200 0.9500 0.9900 1.0200 ;
    END
    ANTENNAGATEAREA 0.1146 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.6500 1.0200 0.7500 ;
        RECT 0.0450 0.7500 0.1450 1.6400 ;
        RECT 0.8500 0.4600 1.0200 0.6500 ;
        RECT 0.3400 0.4150 0.4300 0.6500 ;
        RECT 0.0450 1.6400 0.9200 1.7400 ;
        RECT 0.7500 1.7400 0.9200 1.9300 ;
    END
    ANTENNADIFFAREA 0.3522 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5250 1.2600 1.2150 1.3500 ;
        RECT 0.5250 1.2500 1.2950 1.2600 ;
        RECT 0.5250 1.2250 0.6150 1.2500 ;
        RECT 1.1250 1.1700 1.2950 1.2500 ;
        RECT 0.4450 1.1350 0.6150 1.2250 ;
    END
    ANTENNAGATEAREA 0.1146 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.1300 1.8300 0.2200 2.0800 ;
        RECT 1.4300 1.8200 1.5200 2.0800 ;
    END
  END VDD
END NOR3_X1P4A_A12TH

MACRO NOR3_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 1.0900 0.3200 1.1900 0.7600 ;
        RECT 1.6100 0.3200 1.7100 0.7600 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6900 1.2400 1.1100 1.3600 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.6100 1.8450 1.7100 2.0800 ;
        RECT 0.1050 1.7700 0.2050 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 1.3300 1.1500 ;
        RECT 0.4600 1.1500 0.5600 1.2600 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.4500 1.5400 1.5500 ;
        RECT 1.4400 1.0650 1.5400 1.4500 ;
        RECT 0.2100 0.9400 0.3100 1.4500 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 1.6500 1.7500 1.7500 ;
        RECT 0.7950 1.7500 0.9650 1.9800 ;
        RECT 1.6500 0.9500 1.7500 1.6500 ;
        RECT 0.8300 0.8500 1.7500 0.9500 ;
        RECT 0.8300 0.4200 0.9300 0.8500 ;
        RECT 1.3500 0.4200 1.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.26025 ;
  END Y
END NOR3_X1P4M_A12TH

MACRO NOR3_X2A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7800 ;
        RECT 0.6150 0.3200 0.7150 0.6950 ;
        RECT 1.1350 0.3200 1.2350 0.6950 ;
        RECT 1.6550 0.3200 1.7550 0.7100 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 1.6000 1.5500 ;
        RECT 0.2500 0.9900 0.3500 1.4500 ;
        RECT 1.5000 0.9900 1.6000 1.4500 ;
    END
    ANTENNAGATEAREA 0.162 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5050 1.2500 1.3500 1.3500 ;
        RECT 0.5050 0.9900 0.6050 1.2500 ;
        RECT 1.2450 0.9900 1.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.162 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7150 1.0500 1.1350 1.1500 ;
    END
    ANTENNAGATEAREA 0.162 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9000 1.9500 1.6500 ;
        RECT 0.8400 1.6500 1.9500 1.7500 ;
        RECT 0.3550 0.8000 1.9500 0.9000 ;
        RECT 0.8400 1.7500 1.0100 1.9600 ;
        RECT 0.3550 0.4250 0.4550 0.8000 ;
        RECT 0.8750 0.4250 0.9750 0.8000 ;
        RECT 1.3950 0.4250 1.4950 0.8000 ;
    END
    ANTENNADIFFAREA 0.446 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.6550 1.8400 1.7550 2.0800 ;
        RECT 0.0950 1.7700 0.1950 2.0800 ;
    END
  END VDD
END NOR3_X2A_A12TH

MACRO NOR3_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 1.0850 0.3200 1.1850 0.5600 ;
        RECT 1.6050 0.3200 1.7050 0.5600 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 1.2950 1.3500 ;
        RECT 1.1950 1.0400 1.2950 1.2500 ;
        RECT 0.4500 0.8000 0.5550 1.2500 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.4500 1.5550 1.5500 ;
        RECT 1.4550 1.0600 1.5550 1.4500 ;
        RECT 0.2100 0.7800 0.3100 1.4500 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.6500 1.7500 1.7500 ;
        RECT 0.7900 1.7500 0.9600 1.9800 ;
        RECT 1.6500 0.7500 1.7500 1.6500 ;
        RECT 0.7900 0.6500 1.7500 0.7500 ;
        RECT 0.7900 0.4600 0.9600 0.6500 ;
    END
    ANTENNADIFFAREA 0.3695 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.6050 1.8450 1.7050 2.0800 ;
        RECT 0.1050 1.7700 0.2050 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6700 1.0400 1.0850 1.1600 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END A
END NOR3_X2M_A12TH

MACRO NOR3_X3A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.3050 0.3200 0.4750 0.5300 ;
        RECT 0.8250 0.3200 0.9950 0.5300 ;
        RECT 1.3450 0.3200 1.5150 0.5300 ;
        RECT 1.8650 0.3200 2.0350 0.5300 ;
        RECT 2.4200 0.3200 2.5200 0.4100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 1.0500 2.3600 1.1500 ;
        RECT 2.2600 0.9400 2.3600 1.0500 ;
    END
    ANTENNAGATEAREA 0.243 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.7500 2.5500 1.2500 ;
        RECT 1.3800 1.2500 2.5500 1.3500 ;
        RECT 0.0800 0.6500 2.5500 0.7500 ;
        RECT 1.3800 1.3500 1.4800 1.7000 ;
        RECT 2.4200 1.3500 2.5500 1.7350 ;
        RECT 0.0800 0.4300 0.1800 0.6500 ;
        RECT 0.6000 0.4300 0.7000 0.6500 ;
        RECT 1.1200 0.4300 1.2200 0.6500 ;
        RECT 1.6400 0.4300 1.7400 0.6500 ;
        RECT 2.1600 0.4300 2.2600 0.6500 ;
    END
    ANTENNADIFFAREA 0.75675 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9600 0.8500 2.1400 0.9500 ;
    END
    ANTENNAGATEAREA 0.243 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.0800 1.7700 0.1800 2.0800 ;
        RECT 0.6000 1.7700 0.7000 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0500 0.7500 1.1500 ;
    END
    ANTENNAGATEAREA 0.243 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.8600 1.8200 2.0000 1.9200 ;
      RECT 1.9000 1.5100 2.0000 1.8200 ;
      RECT 0.3400 1.4500 0.9600 1.5500 ;
      RECT 0.8600 1.5500 0.9600 1.8200 ;
      RECT 0.3400 1.5500 0.4400 1.8800 ;
  END
END NOR3_X3A_A12TH

MACRO NOR3_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 1.4500 0.3200 1.5400 0.5800 ;
        RECT 1.9700 0.3200 2.0600 0.5800 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3050 1.0500 1.6750 1.1500 ;
        RECT 1.3050 0.7600 1.3950 1.0500 ;
        RECT 0.1850 0.6700 1.3950 0.7600 ;
        RECT 0.1850 0.7600 0.2750 0.8800 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.2100 2.1500 1.4200 ;
        RECT 0.8700 1.4200 2.1500 1.5100 ;
        RECT 2.0600 1.0500 2.1500 1.2100 ;
        RECT 0.8700 1.1800 0.9600 1.4200 ;
        RECT 0.5750 1.0900 0.9600 1.1800 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9400 1.1500 1.2400 ;
        RECT 1.0500 1.2400 1.9050 1.3300 ;
        RECT 0.6050 0.8500 1.1500 0.9400 ;
        RECT 1.8150 1.0500 1.9050 1.2400 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7750 1.6500 2.3550 1.7500 ;
        RECT 0.7750 1.7500 0.8650 1.9900 ;
        RECT 2.1750 1.7500 2.3200 1.9700 ;
        RECT 0.7750 1.6200 0.8650 1.6500 ;
        RECT 2.1750 1.6000 2.3550 1.6500 ;
        RECT 2.2650 0.9600 2.3550 1.6000 ;
        RECT 1.7100 0.8700 2.3550 0.9600 ;
        RECT 2.2300 0.5900 2.3200 0.8700 ;
        RECT 1.7100 0.5800 1.8000 0.8700 ;
    END
    ANTENNADIFFAREA 0.5976 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0800 1.8400 0.1700 2.0800 ;
        RECT 1.4500 1.8400 1.5400 2.0800 ;
    END
  END VDD
END NOR3_X3M_A12TH

MACRO NOR3_X4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.6300 ;
        RECT 0.5650 0.3200 0.7350 0.5300 ;
        RECT 1.0850 0.3200 1.2550 0.5300 ;
        RECT 1.6050 0.3200 1.7750 0.5300 ;
        RECT 2.1250 0.3200 2.2950 0.5300 ;
        RECT 2.6450 0.3200 2.8150 0.5300 ;
        RECT 3.2000 0.3200 3.3000 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.7500 3.3500 1.2500 ;
        RECT 1.6400 1.2500 3.3500 1.3500 ;
        RECT 0.3400 0.6500 3.3500 0.7500 ;
        RECT 1.6400 1.3500 1.7400 1.7000 ;
        RECT 2.6800 1.3500 2.7800 1.7000 ;
        RECT 0.3400 0.4300 0.4400 0.6500 ;
        RECT 0.8600 0.4300 0.9600 0.6500 ;
        RECT 1.3800 0.4300 1.4800 0.6500 ;
        RECT 1.9000 0.4300 2.0000 0.6500 ;
        RECT 2.4200 0.4300 2.5200 0.6500 ;
        RECT 2.9400 0.4300 3.0400 0.6500 ;
    END
    ANTENNADIFFAREA 0.892 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2300 0.8500 3.1300 0.9500 ;
        RECT 3.0300 0.9500 3.1300 1.1400 ;
    END
    ANTENNAGATEAREA 0.324 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 1.0100 1.1500 ;
    END
    ANTENNAGATEAREA 0.324 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.3400 1.7700 0.4400 2.0800 ;
        RECT 0.8600 1.7700 0.9600 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5000 1.0500 2.9200 1.1500 ;
    END
    ANTENNAGATEAREA 0.324 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.1200 1.8200 3.3000 1.9200 ;
      RECT 3.2000 1.4900 3.3000 1.8200 ;
      RECT 0.0800 1.4550 1.2200 1.5550 ;
      RECT 1.1200 1.5550 1.2200 1.8200 ;
      RECT 2.1600 1.4900 2.2600 1.8200 ;
      RECT 0.0800 1.5550 0.1800 1.8800 ;
      RECT 0.6000 1.5550 0.7000 1.8850 ;
  END
END NOR3_X4A_A12TH

MACRO NOR3_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.9500 0.3200 1.0400 0.6150 ;
        RECT 1.4700 0.3200 1.5600 0.6150 ;
        RECT 1.9900 0.3200 2.0800 0.6150 ;
        RECT 2.5100 0.3200 2.6000 0.6150 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4050 1.0650 1.6950 1.1550 ;
        RECT 0.4050 1.0500 0.7750 1.0650 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 0.8850 1.9250 0.9500 ;
        RECT 0.9350 0.9500 1.9250 0.9750 ;
        RECT 0.4150 0.8250 1.0250 0.8850 ;
        RECT 1.8350 0.9750 1.9250 1.0950 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3250 1.0500 2.7850 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5500 1.2500 2.1050 1.3400 ;
        RECT 0.5500 1.3400 1.5600 1.3500 ;
        RECT 2.0150 0.7950 2.1050 1.2500 ;
        RECT 0.5500 1.3500 0.6400 1.6350 ;
        RECT 1.4700 1.3500 1.5600 1.6350 ;
        RECT 1.2100 0.7050 2.3400 0.7950 ;
        RECT 1.2100 0.4100 1.3000 0.7050 ;
        RECT 1.7300 0.4100 1.8200 0.7050 ;
        RECT 2.2500 0.4100 2.3400 0.7050 ;
    END
    ANTENNADIFFAREA 0.664 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.2500 1.8400 2.3400 2.0800 ;
        RECT 2.7700 1.8400 2.8600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.7250 2.0800 1.8150 ;
      RECT 1.9900 1.5350 2.0800 1.7250 ;
      RECT 1.9900 1.4450 3.1200 1.5350 ;
      RECT 2.5100 1.5350 2.6000 1.8150 ;
      RECT 3.0300 1.5350 3.1200 1.8150 ;
      RECT 0.0800 1.4450 0.1700 1.7250 ;
      RECT 1.0100 1.4450 1.1000 1.7250 ;
  END
END NOR3_X4M_A12TH

MACRO OA211_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.5900 ;
        RECT 1.3250 0.3200 1.4150 0.7900 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0000 1.5500 1.9000 ;
        RECT 1.4500 0.9000 1.6800 1.0000 ;
        RECT 1.5800 0.4300 1.6800 0.9000 ;
    END
    ANTENNADIFFAREA 0.1304 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9700 0.7600 1.3900 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9550 0.1600 1.3500 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9650 0.5500 1.3650 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8100 0.9500 1.0650 ;
        RECT 0.8500 1.0650 1.0850 1.1550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END C0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.5400 1.7350 0.6300 2.0800 ;
        RECT 1.1650 1.7350 1.2550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7550 0.6900 0.8450 ;
      RECT 0.6000 0.4300 0.6900 0.7550 ;
      RECT 0.0800 0.4300 0.1700 0.7550 ;
      RECT 0.0800 1.5000 1.2850 1.5900 ;
      RECT 1.1950 0.9700 1.2850 1.5000 ;
      RECT 1.0750 0.8800 1.2850 0.9700 ;
      RECT 1.0750 0.4300 1.1650 0.8800 ;
      RECT 0.8600 1.5900 0.9500 1.9200 ;
      RECT 0.0800 1.5900 0.1700 1.9100 ;
  END
END OA211_X0P5M_A12TH

MACRO OA211_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6450 ;
        RECT 1.3250 0.3200 1.4150 0.7650 ;
    END
  END VSS

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8100 0.9500 1.0500 ;
        RECT 0.8500 1.0500 1.0850 1.1500 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0000 1.5500 1.7450 ;
        RECT 1.4500 0.9000 1.6800 1.0000 ;
        RECT 1.5800 0.4550 1.6800 0.9000 ;
    END
    ANTENNADIFFAREA 0.1848 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9400 0.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9550 0.1600 1.3500 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.9850 0.7600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.5650 1.7650 0.6650 2.0800 ;
        RECT 1.1550 1.7650 1.2550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7550 0.6900 0.8450 ;
      RECT 0.6000 0.4300 0.6900 0.7550 ;
      RECT 0.0800 0.4300 0.1700 0.7550 ;
      RECT 0.0800 1.5000 1.2850 1.5900 ;
      RECT 1.1950 0.9600 1.2850 1.5000 ;
      RECT 1.0750 0.8700 1.2850 0.9600 ;
      RECT 1.0750 0.4300 1.1650 0.8700 ;
      RECT 0.8600 1.5900 0.9500 1.8850 ;
      RECT 0.0800 1.5900 0.1700 1.9100 ;
  END
END OA211_X0P7M_A12TH

MACRO OA211_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6300 ;
        RECT 1.3250 0.3200 1.4150 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.5350 1.7900 0.6350 2.0800 ;
        RECT 1.1600 1.7900 1.2600 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9850 0.7500 1.2500 ;
        RECT 0.6500 1.2500 0.8500 1.3500 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9550 0.1600 1.3450 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0000 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8100 0.9500 1.0450 ;
        RECT 0.8500 1.0450 1.1350 1.1350 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9100 1.5500 1.8800 ;
        RECT 1.4500 0.8100 1.6800 0.9100 ;
        RECT 1.5800 0.4900 1.6800 0.8100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7550 0.6900 0.8450 ;
      RECT 0.6000 0.4350 0.6900 0.7550 ;
      RECT 0.0800 0.4350 0.1700 0.7550 ;
      RECT 0.0800 1.5000 1.3400 1.5900 ;
      RECT 1.2500 0.9000 1.3400 1.5000 ;
      RECT 1.0750 0.8100 1.3400 0.9000 ;
      RECT 0.0800 1.5900 0.1700 1.9100 ;
      RECT 1.0750 0.4750 1.1650 0.8100 ;
      RECT 0.8550 1.5900 0.9550 1.9650 ;
  END
END OA211_X1M_A12TH

MACRO OA211_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.7350 ;
        RECT 0.8600 0.3200 0.9500 0.7500 ;
        RECT 2.3100 0.3200 2.4000 0.8250 ;
        RECT 2.8300 0.3200 2.9200 0.7600 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.2500 1.0600 1.3500 ;
        RECT 0.9600 1.0550 1.0600 1.2500 ;
    END
    ANTENNAGATEAREA 0.1404 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4050 1.0450 0.8400 1.1550 ;
    END
    ANTENNAGATEAREA 0.1404 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2000 1.2500 2.0400 1.3500 ;
        RECT 1.2000 1.0550 1.3000 1.2500 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 1.0450 1.9300 1.1550 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9500 2.9500 1.2500 ;
        RECT 2.5650 1.2500 2.9500 1.3500 ;
        RECT 2.5650 0.8500 2.9500 0.9500 ;
        RECT 2.5650 1.3500 2.6650 1.8000 ;
        RECT 2.5650 0.4750 2.6650 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.5450 1.6650 0.6350 2.0800 ;
        RECT 1.2650 1.6600 1.3550 2.0800 ;
        RECT 1.7850 1.6600 1.8750 2.0800 ;
        RECT 2.3100 1.5850 2.4000 2.0800 ;
        RECT 2.8300 1.5850 2.9200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8550 1.2100 0.9450 ;
      RECT 1.1200 0.5700 1.2100 0.8550 ;
      RECT 1.1200 0.4800 2.2100 0.5700 ;
      RECT 0.0800 0.4150 0.1700 0.8550 ;
      RECT 0.6000 0.4150 0.6900 0.8550 ;
      RECT 2.1300 1.0600 2.7400 1.1500 ;
      RECT 0.0800 1.5700 0.1700 1.8900 ;
      RECT 1.0050 1.5700 1.0950 1.7550 ;
      RECT 1.5250 1.5700 1.6150 1.7550 ;
      RECT 0.0800 1.4800 2.2200 1.5700 ;
      RECT 2.0600 1.5700 2.1500 1.7550 ;
      RECT 2.1300 1.1500 2.2200 1.4800 ;
      RECT 2.1300 0.7700 2.2200 1.0600 ;
      RECT 1.5200 0.6800 2.2200 0.7700 ;
  END
END OA211_X1P4M_A12TH

MACRO OA211_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6200 ;
        RECT 0.8600 0.3200 0.9500 0.6200 ;
        RECT 2.3650 0.3200 2.4550 0.6450 ;
        RECT 2.8850 0.3200 2.9750 0.6450 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9500 2.9500 1.2500 ;
        RECT 2.6150 1.2500 2.9500 1.3500 ;
        RECT 2.6200 0.8500 2.9500 0.9500 ;
        RECT 2.6150 1.3500 2.7150 1.7400 ;
        RECT 2.6200 0.4950 2.7200 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3950 1.2500 1.8150 1.3500 ;
    END
    ANTENNAGATEAREA 0.1326 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1550 1.0500 2.0400 1.1500 ;
        RECT 1.9400 1.1500 2.0400 1.2650 ;
    END
    ANTENNAGATEAREA 0.1326 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.1800 0.8250 1.3500 ;
    END
    ANTENNAGATEAREA 0.1842 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0250 0.3550 1.3050 ;
        RECT 0.2450 0.9150 1.0650 1.0250 ;
        RECT 0.9550 1.0250 1.0650 1.2500 ;
    END
    ANTENNAGATEAREA 0.1842 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.3650 1.7700 2.4550 2.0800 ;
        RECT 2.8850 1.7700 2.9750 2.0800 ;
        RECT 0.6000 1.7650 0.6900 2.0800 ;
        RECT 1.3200 1.6750 1.4100 2.0800 ;
        RECT 1.8400 1.6750 1.9300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7150 1.2100 0.8050 ;
      RECT 1.1200 0.5700 1.2100 0.7150 ;
      RECT 1.1200 0.4800 2.1950 0.5700 ;
      RECT 0.0800 0.4150 0.1700 0.7150 ;
      RECT 0.6000 0.4150 0.6900 0.7150 ;
      RECT 2.1350 1.0600 2.6650 1.1500 ;
      RECT 0.1350 1.5850 0.2250 1.9250 ;
      RECT 1.0600 1.5850 1.1500 1.9100 ;
      RECT 1.5800 1.5850 1.6700 1.9100 ;
      RECT 0.1350 1.4950 2.2250 1.5850 ;
      RECT 2.1000 1.5850 2.1900 1.9100 ;
      RECT 2.1350 1.1500 2.2250 1.4950 ;
      RECT 2.1350 0.7700 2.2250 1.0600 ;
      RECT 1.5200 0.6800 2.2250 0.7700 ;
  END
END OA211_X2M_A12TH

MACRO OA211_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.5900 ;
        RECT 0.8600 0.3200 0.9500 0.5900 ;
        RECT 1.3800 0.3200 1.4700 0.5900 ;
        RECT 3.3700 0.3200 3.4600 0.6200 ;
        RECT 3.9150 0.3200 4.0050 0.6200 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.2500 1.5800 1.3500 ;
        RECT 0.7000 1.1850 0.8000 1.2500 ;
        RECT 1.4800 1.0800 1.5800 1.2500 ;
        RECT 0.5350 1.0850 0.8000 1.1850 ;
    END
    ANTENNAGATEAREA 0.2799 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1450 1.1000 0.3500 1.1900 ;
        RECT 0.2500 0.9700 0.3500 1.1000 ;
        RECT 0.2500 0.8700 1.0300 0.9700 ;
        RECT 0.9300 0.9700 1.0300 1.0550 ;
        RECT 0.9300 1.0550 1.3500 1.1550 ;
    END
    ANTENNAGATEAREA 0.2799 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7250 1.4500 2.8450 1.5500 ;
        RECT 1.7250 1.1100 1.8250 1.4500 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9450 1.0500 3.0800 1.1500 ;
        RECT 2.9800 1.1500 3.0800 1.4900 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9300 4.3500 1.2500 ;
        RECT 3.6500 1.2500 4.3500 1.3500 ;
        RECT 3.6500 0.8300 4.3500 0.9300 ;
        RECT 3.6500 1.3500 3.7500 1.7400 ;
        RECT 4.1750 1.3500 4.2650 1.7400 ;
        RECT 4.1750 0.4950 4.2650 0.8300 ;
        RECT 3.6500 0.4850 3.7500 0.8300 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 1.8400 1.8800 1.9300 2.0800 ;
        RECT 2.3600 1.8800 2.4500 2.0800 ;
        RECT 2.8800 1.8800 2.9700 2.0800 ;
        RECT 1.1200 1.8400 1.2100 2.0800 ;
        RECT 3.3950 1.7700 3.4850 2.0800 ;
        RECT 3.9150 1.7700 4.0050 2.0800 ;
        RECT 0.1400 1.7650 0.2300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6900 1.7300 0.7800 ;
      RECT 1.6400 0.5750 1.7300 0.6900 ;
      RECT 1.6400 0.4850 2.7100 0.5750 ;
      RECT 0.0800 0.4100 0.1700 0.6900 ;
      RECT 0.6000 0.4100 0.6900 0.6900 ;
      RECT 1.1200 0.4100 1.2100 0.6900 ;
      RECT 3.2000 1.0600 3.9650 1.1500 ;
      RECT 1.5800 1.7500 1.6700 1.9150 ;
      RECT 2.1000 1.7500 2.1900 1.9150 ;
      RECT 2.6200 1.7500 2.7100 1.9150 ;
      RECT 0.5600 1.6600 3.2900 1.7500 ;
      RECT 3.1400 1.7500 3.2300 1.9150 ;
      RECT 3.2000 1.1500 3.2900 1.6600 ;
      RECT 3.2000 0.8400 3.2900 1.0600 ;
      RECT 2.0350 0.7500 3.2900 0.8400 ;
      RECT 3.0200 0.4700 3.1100 0.7500 ;
      RECT 0.5600 1.4600 0.7300 1.6600 ;
  END
END OA211_X3M_A12TH

MACRO OA211_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3450 0.3200 0.4350 0.6100 ;
        RECT 0.8650 0.3200 0.9550 0.6100 ;
        RECT 1.3850 0.3200 1.4750 0.6100 ;
        RECT 1.9050 0.3200 1.9950 0.6100 ;
        RECT 4.3600 0.3200 4.4500 0.6400 ;
        RECT 4.9050 0.3200 4.9950 0.6400 ;
        RECT 5.4250 0.3200 5.5150 0.6400 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.9850 0.3500 1.2300 ;
        RECT 0.2450 0.8850 2.1000 0.9850 ;
        RECT 1.0100 0.9850 1.2200 1.1500 ;
        RECT 2.0000 0.9850 2.1000 1.3000 ;
    END
    ANTENNAGATEAREA 0.3708 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.2500 1.5400 1.3500 ;
        RECT 0.7050 1.2150 0.8050 1.2500 ;
        RECT 1.4400 1.2000 1.5400 1.2500 ;
        RECT 0.5150 1.1150 0.8050 1.2150 ;
        RECT 1.4400 1.1100 1.8100 1.2000 ;
    END
    ANTENNAGATEAREA 0.3708 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5450 1.0500 3.5300 1.1500 ;
        RECT 3.4300 1.1500 3.5300 1.2500 ;
        RECT 3.4300 1.2500 3.8400 1.3500 ;
    END
    ANTENNAGATEAREA 0.2664 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2200 1.4500 4.1250 1.5500 ;
        RECT 2.2200 1.3550 2.3200 1.4500 ;
        RECT 4.0250 1.0200 4.1250 1.4500 ;
    END
    ANTENNAGATEAREA 0.2664 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 0.9500 5.3500 1.2500 ;
        RECT 4.6400 1.2500 5.3500 1.3500 ;
        RECT 4.6400 0.8500 5.3500 0.9500 ;
        RECT 4.6400 1.3500 4.7400 1.7200 ;
        RECT 5.1650 1.3500 5.2550 1.7200 ;
        RECT 4.6400 0.4950 4.7400 0.8500 ;
        RECT 5.1650 0.4950 5.2550 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 2.3100 1.8600 2.4000 2.0800 ;
        RECT 2.8350 1.8600 2.9250 2.0800 ;
        RECT 3.3550 1.8600 3.4450 2.0800 ;
        RECT 3.8750 1.8600 3.9650 2.0800 ;
        RECT 4.3850 1.8250 4.4750 2.0800 ;
        RECT 0.6050 1.7700 0.6950 2.0800 ;
        RECT 1.5750 1.7700 1.6650 2.0800 ;
        RECT 4.9050 1.7700 4.9950 2.0800 ;
        RECT 5.4250 1.7700 5.5150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0850 0.7000 2.2550 0.7900 ;
      RECT 2.1650 0.5700 2.2550 0.7000 ;
      RECT 2.1650 0.4800 4.1650 0.5700 ;
      RECT 0.0850 0.4100 0.1750 0.7000 ;
      RECT 0.6050 0.4100 0.6950 0.7000 ;
      RECT 1.1250 0.4100 1.2150 0.7000 ;
      RECT 1.6450 0.4100 1.7350 0.7000 ;
      RECT 4.2750 1.0550 5.1400 1.1450 ;
      RECT 0.1450 1.5850 0.2350 1.9300 ;
      RECT 1.0850 1.5850 1.1750 1.9300 ;
      RECT 2.0450 1.7300 2.1350 1.9100 ;
      RECT 1.8150 1.5850 1.9050 1.6400 ;
      RECT 0.1450 1.4950 1.9050 1.5850 ;
      RECT 2.5750 1.7300 2.6650 1.9100 ;
      RECT 3.0950 1.7300 3.1850 1.9100 ;
      RECT 3.6150 1.7300 3.7050 1.9100 ;
      RECT 1.8150 1.6400 4.3650 1.7300 ;
      RECT 4.1350 1.7300 4.2250 1.9100 ;
      RECT 4.2750 1.1450 4.3650 1.6400 ;
      RECT 4.2750 0.8350 4.3650 1.0550 ;
      RECT 2.5600 0.7450 4.3650 0.8350 ;
  END
END OA211_X4M_A12TH

MACRO OA211_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.3450 0.3200 0.4350 0.5800 ;
        RECT 0.8650 0.3200 0.9550 0.5800 ;
        RECT 1.3850 0.3200 1.4750 0.5800 ;
        RECT 1.9050 0.3200 1.9950 0.5800 ;
        RECT 2.4250 0.3200 2.5150 0.5800 ;
        RECT 2.9450 0.3200 3.0350 0.5800 ;
        RECT 6.4500 0.3200 6.5400 0.6500 ;
        RECT 6.9900 0.3200 7.0800 0.6400 ;
        RECT 7.5100 0.3200 7.6000 0.6400 ;
        RECT 8.0300 0.3200 8.1200 0.6400 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 1.0500 1.9000 1.1500 ;
        RECT 1.4400 1.1500 1.5500 1.2500 ;
        RECT 1.8000 1.1500 1.9000 1.2500 ;
        RECT 0.8500 1.2500 1.5500 1.3500 ;
        RECT 1.8000 1.2500 2.7100 1.3500 ;
        RECT 0.8500 1.1500 0.9500 1.2500 ;
        RECT 2.6100 1.2400 2.7100 1.2500 ;
        RECT 0.4950 1.0500 0.9500 1.1500 ;
        RECT 2.6100 1.1400 2.8250 1.2400 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1300 1.0800 0.3500 1.1900 ;
        RECT 0.2450 0.9500 0.3500 1.0800 ;
        RECT 0.2450 0.8500 2.1100 0.9500 ;
        RECT 1.0900 0.9500 1.2600 1.1500 ;
        RECT 2.0100 0.9500 2.1100 1.0500 ;
        RECT 2.0100 1.0500 2.5000 1.1500 ;
        RECT 2.4000 0.9500 2.5000 1.0500 ;
        RECT 2.4000 0.8500 3.1150 0.9500 ;
        RECT 3.0150 0.9500 3.1150 1.3550 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2600 1.2500 6.1950 1.3500 ;
        RECT 3.2600 1.3500 3.3600 1.5600 ;
    END
    ANTENNAGATEAREA 0.3996 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5250 1.0500 5.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.3996 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8500 0.9500 7.9500 1.2500 ;
        RECT 6.7250 1.2500 7.9500 1.3500 ;
        RECT 6.7250 0.8500 7.9500 0.9500 ;
        RECT 6.7250 1.3500 6.8250 1.7550 ;
        RECT 7.2500 1.3500 7.3400 1.7200 ;
        RECT 7.7700 1.3500 7.8600 1.7200 ;
        RECT 6.7250 0.5050 6.8250 0.8500 ;
        RECT 7.2500 0.4850 7.3400 0.8500 ;
        RECT 7.7700 0.4850 7.8600 0.8500 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 3.3600 1.8750 3.4500 2.0800 ;
        RECT 3.8800 1.8750 3.9700 2.0800 ;
        RECT 4.4000 1.8750 4.4900 2.0800 ;
        RECT 4.9200 1.8750 5.0100 2.0800 ;
        RECT 5.4400 1.8750 5.5300 2.0800 ;
        RECT 5.9600 1.8750 6.0500 2.0800 ;
        RECT 6.4700 1.8150 6.5600 2.0800 ;
        RECT 0.6050 1.7700 0.6950 2.0800 ;
        RECT 1.6450 1.7700 1.7350 2.0800 ;
        RECT 2.6250 1.7700 2.7150 2.0800 ;
        RECT 6.9900 1.7700 7.0800 2.0800 ;
        RECT 7.5100 1.7700 7.6000 2.0800 ;
        RECT 8.0300 1.7700 8.1200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0850 0.6700 3.3000 0.7600 ;
      RECT 3.2100 0.5850 3.3000 0.6700 ;
      RECT 3.2100 0.4950 6.2900 0.5850 ;
      RECT 0.0850 0.4850 0.1750 0.6700 ;
      RECT 0.5650 0.4100 0.7350 0.6700 ;
      RECT 1.0850 0.4100 1.2550 0.6700 ;
      RECT 1.6050 0.4100 1.7750 0.6700 ;
      RECT 2.1250 0.4100 2.2950 0.6700 ;
      RECT 2.6450 0.4100 2.8150 0.6700 ;
      RECT 6.3100 1.0700 7.7100 1.1600 ;
      RECT 3.1000 1.7500 3.1900 1.9150 ;
      RECT 2.9850 1.6450 3.0750 1.6600 ;
      RECT 1.1250 1.5550 3.0750 1.6450 ;
      RECT 3.6200 1.7500 3.7100 1.9150 ;
      RECT 4.1400 1.7500 4.2300 1.9150 ;
      RECT 4.6600 1.7500 4.7500 1.9150 ;
      RECT 5.1800 1.7500 5.2700 1.9150 ;
      RECT 5.7000 1.7500 5.7900 1.9150 ;
      RECT 2.9850 1.6600 6.4000 1.7500 ;
      RECT 6.2200 1.7500 6.3100 1.9150 ;
      RECT 6.3100 1.1600 6.4000 1.6600 ;
      RECT 6.3100 0.8400 6.4000 1.0700 ;
      RECT 3.6100 0.7500 6.4000 0.8400 ;
      RECT 0.1450 1.5450 0.2350 1.8850 ;
      RECT 1.1250 1.6450 1.2150 1.8850 ;
      RECT 1.1250 1.5450 1.2150 1.5550 ;
      RECT 0.1450 1.4550 1.2150 1.5450 ;
      RECT 2.1650 1.6450 2.2550 1.9600 ;
  END
END OA211_X6M_A12TH

MACRO OA21_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.9100 0.3200 1.0000 0.6900 ;
        RECT 0.3550 0.3200 0.4450 0.5950 ;
        RECT 0.9100 0.6900 1.1200 0.7800 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.2300 1.6400 1.3200 2.0800 ;
        RECT 0.3650 1.5300 0.5750 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6200 1.2550 ;
        RECT 0.5300 0.9050 0.6200 1.0100 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7300 1.0500 1.0550 1.1500 ;
        RECT 0.8150 1.1500 0.9050 1.2600 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2450 1.2750 1.3500 1.5100 ;
        RECT 1.1650 1.1650 1.3500 1.2750 ;
        RECT 1.1650 1.0700 1.2550 1.1650 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5350 0.1500 1.7650 ;
        RECT 0.0500 1.7650 0.1700 1.9550 ;
        RECT 0.0500 0.4450 0.2450 0.5350 ;
    END
    ANTENNADIFFAREA 0.1358 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7100 1.4400 0.8000 1.8300 ;
      RECT 0.2400 1.3500 0.8000 1.4400 ;
      RECT 0.2400 0.7050 0.6000 0.7950 ;
      RECT 0.2400 0.7950 0.3300 1.3500 ;
      RECT 0.7100 0.8700 1.3200 0.9600 ;
      RECT 1.2300 0.7500 1.3200 0.8700 ;
      RECT 0.7100 0.7500 0.8000 0.8700 ;
  END
END OA21_X0P5M_A12TH

MACRO OA21_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4600 0.4850 ;
        RECT 1.1400 0.3200 1.2600 0.7700 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.7900 1.3050 ;
    END
    ANTENNAGATEAREA 0.0405 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0900 0.5500 1.5100 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.4500 1.5500 1.9050 ;
        RECT 1.4100 0.4450 1.5200 1.4500 ;
    END
    ANTENNADIFFAREA 0.202125 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 0.8100 0.3500 0.9200 ;
        RECT 0.2400 0.9200 0.3500 1.1200 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8700 1.8850 0.9700 2.0800 ;
        RECT 1.1500 1.7000 1.2500 2.0800 ;
        RECT 0.0900 1.6800 0.1900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 0.5950 0.7050 0.6950 ;
      RECT 0.6150 0.4400 0.7050 0.5950 ;
      RECT 0.0950 0.4400 0.1850 0.5950 ;
      RECT 0.9200 1.0450 1.3000 1.1450 ;
      RECT 0.5700 1.7850 0.6600 1.9800 ;
      RECT 0.5700 1.6850 1.0100 1.7850 ;
      RECT 0.9200 1.1450 1.0100 1.6850 ;
      RECT 0.9200 0.5650 1.0100 1.0450 ;
      RECT 0.8150 0.4750 1.0100 0.5650 ;
  END
END OA21_X0P7M_A12TH

MACRO OA21_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4600 0.4300 ;
        RECT 1.1400 0.3200 1.2600 0.6700 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7150 0.7900 1.1150 ;
    END
    ANTENNAGATEAREA 0.0525 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2950 1.2400 0.7050 1.3500 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.2500 1.5500 1.7200 ;
        RECT 1.4100 0.5250 1.5200 1.2500 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.7150 0.3500 1.1150 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8700 1.9900 0.9700 2.0800 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 1.1500 1.7700 1.2500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 0.5350 0.7050 0.6250 ;
      RECT 0.6150 0.4150 0.7050 0.5350 ;
      RECT 0.0950 0.4150 0.1850 0.5350 ;
      RECT 0.9350 1.0750 1.3000 1.1750 ;
      RECT 0.5700 1.7900 0.6600 1.9900 ;
      RECT 0.5700 1.7000 1.0250 1.7900 ;
      RECT 0.9350 1.1750 1.0250 1.7000 ;
      RECT 0.9350 0.5650 1.0250 1.0750 ;
      RECT 0.8150 0.4750 1.0250 0.5650 ;
  END
END OA21_X1M_A12TH

MACRO OA21_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.8650 0.3200 1.0350 0.5400 ;
        RECT 1.4700 0.3200 1.5600 0.8900 ;
        RECT 1.9900 0.3200 2.0800 0.8400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7300 1.4500 2.1550 1.5500 ;
        RECT 1.7300 1.5500 1.8200 1.9300 ;
        RECT 2.0650 1.0450 2.1550 1.4500 ;
        RECT 1.7700 0.9550 2.1550 1.0450 ;
        RECT 1.6900 0.6650 1.8600 0.9550 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.0500 1.3600 1.1500 ;
        RECT 1.2700 1.1500 1.3600 1.1800 ;
        RECT 1.2700 0.9700 1.3600 1.0500 ;
    END
    ANTENNAGATEAREA 0.1068 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9300 0.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.2500 1.1300 1.3500 ;
    END
    ANTENNAGATEAREA 0.1068 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.9900 1.7150 2.0800 2.0800 ;
        RECT 1.4700 1.6600 1.5600 2.0800 ;
        RECT 0.3550 1.6500 0.4450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 0.6300 1.2950 0.7200 ;
      RECT 1.1250 0.7200 1.2950 0.7700 ;
      RECT 1.1250 0.4800 1.2950 0.6300 ;
      RECT 0.3550 0.7200 0.4450 0.8400 ;
      RECT 0.6450 0.7200 0.7350 0.8100 ;
      RECT 0.3550 0.4700 0.4450 0.6300 ;
      RECT 0.6450 0.4400 0.7350 0.6300 ;
      RECT 1.5500 1.2700 1.9550 1.3600 ;
      RECT 0.0500 1.4400 1.6400 1.5300 ;
      RECT 1.5500 1.3600 1.6400 1.4400 ;
      RECT 0.0950 1.5800 0.1850 1.9300 ;
      RECT 0.0500 1.5300 0.1850 1.5800 ;
      RECT 0.0500 0.8400 0.1400 1.4400 ;
      RECT 0.0500 0.7500 0.1850 0.8400 ;
      RECT 0.0950 0.4500 0.1850 0.7500 ;
      RECT 0.9050 1.5300 0.9950 1.9300 ;
  END
END OA21_X1P4M_A12TH

MACRO OA21_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.5650 ;
        RECT 0.8600 0.3200 0.9500 0.5650 ;
        RECT 1.9050 0.3200 1.9950 0.6700 ;
        RECT 2.4250 0.3200 2.5150 0.6700 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.2500 0.8900 1.3600 ;
    END
    ANTENNAGATEAREA 0.1404 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8900 1.5500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0996 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9400 2.3500 1.4500 ;
        RECT 2.1600 1.4500 2.3500 1.5500 ;
        RECT 2.1600 0.8400 2.3500 0.9400 ;
        RECT 2.1600 1.5500 2.2600 1.8800 ;
        RECT 2.1600 0.5100 2.2600 0.8400 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.0350 0.3800 1.1900 ;
        RECT 0.2250 0.9450 1.0600 1.0350 ;
        RECT 0.9600 1.0350 1.0600 1.1150 ;
    END
    ANTENNAGATEAREA 0.1404 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 1.1200 1.7800 1.2100 2.0800 ;
        RECT 1.6400 1.7800 1.7300 2.0800 ;
        RECT 1.9050 1.7700 1.9950 2.0800 ;
        RECT 2.4250 1.7700 2.5150 2.0800 ;
        RECT 0.0800 1.7350 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7200 1.2100 0.8200 ;
      RECT 1.1200 0.5700 1.2100 0.7200 ;
      RECT 1.1200 0.4800 1.7900 0.5700 ;
      RECT 0.0800 0.4100 0.1700 0.7200 ;
      RECT 0.6000 0.4100 0.6900 0.7200 ;
      RECT 1.6900 1.0750 2.1400 1.1650 ;
      RECT 0.6000 1.6500 0.6900 1.9900 ;
      RECT 1.3800 1.6500 1.4700 1.9900 ;
      RECT 0.6000 1.5600 1.7800 1.6500 ;
      RECT 1.6900 1.1650 1.7800 1.5600 ;
      RECT 1.6900 0.7750 1.7800 1.0750 ;
      RECT 1.3200 0.6850 1.7800 0.7750 ;
  END
END OA21_X2M_A12TH

MACRO OA21_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.8600 0.3200 0.9500 0.6250 ;
        RECT 1.1950 0.3200 1.2850 0.6000 ;
        RECT 1.7150 0.3200 1.8050 0.6000 ;
        RECT 2.2500 0.3200 2.3400 0.6750 ;
        RECT 2.7700 0.3200 2.8600 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.7700 1.7700 2.8600 2.0800 ;
        RECT 1.7150 1.6900 1.8050 2.0800 ;
        RECT 2.2500 1.6200 2.3400 2.0800 ;
        RECT 0.3400 1.4900 0.4300 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0500 0.7900 1.1950 ;
    END
    ANTENNAGATEAREA 0.1518 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9050 1.0500 1.3300 1.1650 ;
    END
    ANTENNAGATEAREA 0.2127 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5700 1.0500 2.0300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2127 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5100 1.2500 3.1200 1.3500 ;
        RECT 2.5100 1.3500 2.6000 1.7200 ;
        RECT 3.0300 1.3500 3.1200 1.7150 ;
        RECT 3.0300 0.9800 3.1200 1.2500 ;
        RECT 2.5100 0.8900 3.1200 0.9800 ;
        RECT 2.5100 0.5300 2.6000 0.8900 ;
        RECT 3.0300 0.5300 3.1200 0.8900 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.4550 1.5100 2.0650 1.6000 ;
      RECT 1.9750 1.6000 2.0650 1.9400 ;
      RECT 0.9350 1.8100 1.5450 1.9000 ;
      RECT 1.4550 1.6000 1.5450 1.8100 ;
      RECT 0.9350 1.4900 1.0250 1.8100 ;
      RECT 0.6000 0.7150 2.0650 0.8050 ;
      RECT 1.9750 0.4350 2.0650 0.7150 ;
      RECT 0.6000 0.5700 0.6900 0.7150 ;
      RECT 0.0800 0.4800 0.6900 0.5700 ;
      RECT 0.0800 0.5700 0.1700 0.6900 ;
      RECT 0.6000 0.4350 0.6900 0.4800 ;
      RECT 1.4550 0.4350 1.5450 0.7150 ;
      RECT 2.3300 1.0700 2.8050 1.1600 ;
      RECT 0.0800 1.3750 0.1700 1.7650 ;
      RECT 0.0800 0.9500 0.1700 1.2850 ;
      RECT 1.1950 1.3750 1.2850 1.6800 ;
      RECT 0.6750 1.3750 0.7650 1.7650 ;
      RECT 0.0800 0.8600 0.4700 0.9500 ;
      RECT 0.3000 0.6600 0.4700 0.8600 ;
      RECT 0.0800 1.2850 2.4200 1.3750 ;
      RECT 2.3300 1.1600 2.4200 1.2850 ;
  END
END OA21_X3M_A12TH

MACRO OA21_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4600 0.5800 ;
        RECT 0.8600 0.3200 0.9800 0.5800 ;
        RECT 1.3800 0.3200 1.5000 0.5800 ;
        RECT 2.7250 0.3200 2.8350 0.6700 ;
        RECT 3.2450 0.3200 3.3550 0.6700 ;
        RECT 3.7650 0.3200 3.8750 0.6700 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8450 0.8900 1.9550 1.3100 ;
    END
    ANTENNAGATEAREA 0.1917 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5500 1.0500 1.6000 1.1600 ;
        RECT 1.4900 0.9250 1.6000 1.0500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9900 0.8500 3.7500 0.9500 ;
        RECT 3.6500 0.9500 3.7500 1.2950 ;
        RECT 2.9900 0.5100 3.0900 0.8500 ;
        RECT 3.5100 0.5100 3.6100 0.8500 ;
        RECT 2.9900 1.2950 3.7500 1.3850 ;
        RECT 2.9900 1.3850 3.0900 1.7250 ;
        RECT 3.5150 1.3850 3.6050 1.7050 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8500 1.2850 0.9600 ;
        RECT 0.2400 0.9600 0.3500 1.1100 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 1.1300 1.9900 1.2300 2.0800 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 1.9300 1.7700 2.0300 2.0800 ;
        RECT 2.4500 1.7700 2.5500 2.0800 ;
        RECT 2.7300 1.7700 2.8300 2.0800 ;
        RECT 3.2500 1.7700 3.3500 2.0800 ;
        RECT 3.7700 1.7700 3.8700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 1.7950 1.5450 1.8850 ;
      RECT 0.3550 1.4950 0.4450 1.7950 ;
      RECT 0.0550 0.6700 1.7450 0.7600 ;
      RECT 1.6550 0.5700 1.7450 0.6700 ;
      RECT 1.6550 0.4800 2.3450 0.5700 ;
      RECT 0.0550 0.4100 0.2250 0.6700 ;
      RECT 0.5750 0.4100 0.7450 0.6700 ;
      RECT 1.0950 0.4100 1.2650 0.6700 ;
      RECT 2.4550 1.0650 3.3250 1.1750 ;
      RECT 1.6550 1.6000 1.7450 1.9500 ;
      RECT 2.1950 1.6000 2.2850 1.9500 ;
      RECT 0.5550 1.5100 2.5450 1.6000 ;
      RECT 2.4550 1.1750 2.5450 1.5100 ;
      RECT 2.4550 0.7900 2.5450 1.0650 ;
      RECT 1.8750 0.6800 2.5450 0.7900 ;
      RECT 2.4550 0.4100 2.5450 0.6800 ;
  END
END OA21_X4M_A12TH

MACRO OA21_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.1500 0.3200 0.2400 0.6850 ;
        RECT 0.6700 0.3200 0.7600 0.6850 ;
        RECT 1.1900 0.3200 1.2800 0.6850 ;
        RECT 1.7100 0.3200 1.8000 0.6850 ;
        RECT 3.2600 0.3200 3.3500 0.5800 ;
        RECT 3.5000 0.3200 3.6700 0.5300 ;
        RECT 4.0600 0.3200 4.1500 0.5800 ;
        RECT 4.5800 0.3200 4.6700 0.5800 ;
        RECT 5.1000 0.3200 5.1900 0.5800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3050 1.4500 1.5400 1.5400 ;
        RECT 0.4100 1.5400 1.5400 1.5500 ;
        RECT 0.3050 0.9800 0.3950 1.4500 ;
        RECT 0.4100 1.5500 0.5000 1.8800 ;
        RECT 0.9300 1.5500 1.0200 1.8800 ;
        RECT 1.4500 1.5500 1.5400 1.8800 ;
        RECT 0.3050 0.8900 1.5400 0.9800 ;
        RECT 0.4100 0.5400 0.5000 0.8900 ;
        RECT 0.9300 0.5400 1.0200 0.8900 ;
        RECT 1.4500 0.5400 1.5400 0.8900 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2950 0.9700 2.7550 1.1500 ;
    END
    ANTENNAGATEAREA 0.2967 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9200 0.8500 3.7250 0.9450 ;
        RECT 2.9200 0.9450 4.7450 0.9500 ;
        RECT 2.9200 0.9500 3.0100 1.1400 ;
        RECT 3.6350 0.9500 4.0450 1.0900 ;
        RECT 4.6550 0.9500 4.7450 0.9900 ;
        RECT 3.9550 0.8500 4.7450 0.9450 ;
        RECT 2.8950 1.1400 3.0100 1.3500 ;
        RECT 4.6550 0.9900 5.0450 1.0900 ;
    END
    ANTENNAGATEAREA 0.4164 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2100 1.2500 5.3000 1.3500 ;
        RECT 3.2100 1.1800 3.6000 1.2500 ;
        RECT 4.1550 1.1800 4.5650 1.2500 ;
        RECT 5.1850 1.0500 5.3000 1.2500 ;
    END
    ANTENNAGATEAREA 0.4164 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.1500 1.7700 0.2400 2.0800 ;
        RECT 0.6700 1.7700 0.7600 2.0800 ;
        RECT 1.1900 1.7700 1.2800 2.0800 ;
        RECT 1.7100 1.7700 1.8000 2.0800 ;
        RECT 3.2800 1.7700 3.3700 2.0800 ;
        RECT 4.3200 1.7700 4.4100 2.0800 ;
        RECT 5.2900 1.7700 5.3800 2.0800 ;
        RECT 2.0100 1.6750 2.1000 2.0800 ;
        RECT 2.5300 1.6750 2.6200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1150 1.4600 4.9200 1.5500 ;
      RECT 4.8300 1.5500 4.9200 1.8900 ;
      RECT 2.2700 1.5500 2.3600 1.8900 ;
      RECT 2.2200 0.6600 2.3100 0.7700 ;
      RECT 2.1150 1.1800 2.2050 1.4600 ;
      RECT 0.4850 1.0900 2.2050 1.1800 ;
      RECT 2.1150 0.8600 2.2050 1.0900 ;
      RECT 2.1150 0.7700 2.8300 0.8600 ;
      RECT 2.7400 0.6600 2.8300 0.7700 ;
      RECT 2.8150 1.5500 2.9050 1.8900 ;
      RECT 3.8000 1.5500 3.8900 1.8900 ;
      RECT 3.0000 0.6700 5.4900 0.7600 ;
      RECT 5.3200 0.4500 5.4900 0.6700 ;
      RECT 1.9600 0.5700 2.0500 0.6800 ;
      RECT 1.9600 0.4800 3.0900 0.5700 ;
      RECT 2.4800 0.5700 2.5700 0.6800 ;
      RECT 3.0000 0.5700 3.0900 0.6700 ;
      RECT 3.7600 0.4500 3.9300 0.6700 ;
      RECT 4.2800 0.4500 4.4500 0.6700 ;
      RECT 4.8000 0.4500 4.9700 0.6700 ;
  END
END OA21_X6M_A12TH

MACRO OA21_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.3750 0.3200 0.4650 0.6150 ;
        RECT 0.8950 0.3200 0.9850 0.6150 ;
        RECT 1.4150 0.3200 1.5050 0.6150 ;
        RECT 1.9350 0.3200 2.0250 0.6150 ;
        RECT 2.4550 0.3200 2.5450 0.6150 ;
        RECT 2.7050 0.3200 2.7950 0.6150 ;
        RECT 4.7250 0.3200 4.8150 0.6750 ;
        RECT 5.2450 0.3200 5.3350 0.6750 ;
        RECT 5.7650 0.3200 5.8550 0.6750 ;
        RECT 6.2850 0.3200 6.3750 0.6750 ;
        RECT 6.8050 0.3200 6.8950 0.6750 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5000 1.0500 0.8700 1.1500 ;
        RECT 0.7800 0.9800 0.8700 1.0500 ;
        RECT 0.7800 0.8900 1.6300 0.9800 ;
        RECT 1.5300 0.9800 1.6300 1.0500 ;
        RECT 1.5300 1.0500 1.9000 1.1500 ;
        RECT 1.8000 0.9800 1.9000 1.0500 ;
        RECT 1.8000 0.8900 2.6100 0.9800 ;
        RECT 2.5200 0.9800 2.6100 1.0600 ;
        RECT 2.5200 1.0600 2.9000 1.1500 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5100 1.0900 4.2300 1.1900 ;
        RECT 3.6100 1.0500 3.7900 1.0900 ;
    END
    ANTENNAGATEAREA 0.3846 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.2500 1.1100 1.3500 ;
        RECT 1.0100 1.2000 1.1100 1.2500 ;
        RECT 0.3000 1.1800 0.3900 1.2500 ;
        RECT 1.0100 1.0700 1.3800 1.2000 ;
        RECT 0.1800 1.0900 0.3900 1.1800 ;
        RECT 1.2800 1.2000 1.3800 1.2500 ;
        RECT 1.2800 1.2500 2.1600 1.3500 ;
        RECT 2.0600 1.1750 2.1600 1.2500 ;
        RECT 2.0600 1.0700 2.4300 1.1750 ;
        RECT 2.3300 1.1750 2.4300 1.2400 ;
        RECT 2.3300 1.2400 3.1000 1.3500 ;
        RECT 3.0100 1.1800 3.1000 1.2400 ;
        RECT 3.0100 1.0900 3.2200 1.1800 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9650 1.2350 6.7650 1.3650 ;
        RECT 4.9650 1.3650 5.0950 1.7200 ;
        RECT 5.4850 1.3650 5.6150 1.7200 ;
        RECT 6.0050 1.3650 6.1350 1.7200 ;
        RECT 6.5250 1.3650 6.6550 1.7200 ;
        RECT 6.6350 0.9650 6.7650 1.2350 ;
        RECT 4.9650 0.8350 6.7650 0.9650 ;
        RECT 4.9650 0.5200 5.0950 0.8350 ;
        RECT 5.4850 0.5200 5.6150 0.8350 ;
        RECT 6.0050 0.5200 6.1350 0.8350 ;
        RECT 6.5250 0.5200 6.6550 0.8350 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 0.1750 1.7700 0.2650 2.0800 ;
        RECT 1.1550 1.7700 1.2450 2.0800 ;
        RECT 2.1950 1.7700 2.2850 2.0800 ;
        RECT 3.1450 1.7700 3.2350 2.0800 ;
        RECT 4.7250 1.7700 4.8150 2.0800 ;
        RECT 5.2450 1.7700 5.3350 2.0800 ;
        RECT 5.7650 1.7700 5.8550 2.0800 ;
        RECT 6.2850 1.7700 6.3750 2.0800 ;
        RECT 6.8050 1.7700 6.8950 2.0800 ;
        RECT 3.6950 1.6550 3.7850 2.0800 ;
        RECT 4.2150 1.6550 4.3050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1150 0.7050 3.1900 0.7950 ;
      RECT 3.0200 0.5700 3.1900 0.7050 ;
      RECT 3.0200 0.4800 4.3450 0.5700 ;
      RECT 3.6550 0.5700 3.8250 0.7700 ;
      RECT 4.1750 0.5700 4.3450 0.7800 ;
      RECT 0.1150 0.4100 0.2050 0.7050 ;
      RECT 0.6350 0.4250 0.7250 0.7050 ;
      RECT 1.1550 0.4250 1.2450 0.7050 ;
      RECT 1.6750 0.4250 1.7650 0.7050 ;
      RECT 2.1950 0.4250 2.2850 0.7050 ;
      RECT 4.4750 1.0550 6.5050 1.1450 ;
      RECT 0.6350 1.5500 0.7250 1.8900 ;
      RECT 1.6750 1.5500 1.7650 1.8900 ;
      RECT 2.6750 1.5500 2.7650 1.8900 ;
      RECT 3.4350 1.5500 3.5250 1.8900 ;
      RECT 3.3950 0.6600 3.5650 0.8700 ;
      RECT 3.9550 1.5500 4.0450 1.8900 ;
      RECT 3.9150 0.6600 4.0850 0.8700 ;
      RECT 0.6350 1.4600 4.5650 1.5500 ;
      RECT 4.4750 1.1450 4.5650 1.4600 ;
      RECT 4.4750 0.9600 4.5650 1.0550 ;
      RECT 3.3950 0.8700 4.5650 0.9600 ;
      RECT 4.4750 0.5350 4.5650 0.8700 ;
  END
END OA21_X8M_A12TH

MACRO OA22_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.7350 ;
        RECT 1.3700 0.3200 1.4600 0.8900 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8900 1.7500 1.4950 ;
        RECT 1.6300 1.4950 1.7500 1.9250 ;
        RECT 1.6300 0.4800 1.7500 0.8900 ;
    END
    ANTENNADIFFAREA 0.1304 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2100 0.1600 1.5950 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.0800 1.7400 0.1700 2.0800 ;
        RECT 1.1200 1.7400 1.2100 2.0800 ;
        RECT 1.3700 1.5200 1.4600 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.2800 1.1800 1.6200 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0400 0.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.2100 0.7650 1.5650 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.0800 0.8300 0.6900 0.9200 ;
      RECT 0.6000 0.5700 0.6900 0.8300 ;
      RECT 0.6000 0.4800 1.2100 0.5700 ;
      RECT 1.1200 0.5700 1.2100 0.7750 ;
      RECT 0.0800 0.6600 0.1700 0.8300 ;
      RECT 0.8600 1.0100 1.5450 1.1000 ;
      RECT 1.4550 1.1000 1.5450 1.4000 ;
      RECT 0.5400 1.8800 0.9500 1.9700 ;
      RECT 0.8600 1.1000 0.9500 1.8800 ;
      RECT 0.8600 0.6900 0.9500 1.0100 ;
  END
END OA22_X0P5M_A12TH

MACRO NOR2_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6950 ;
        RECT 0.6150 0.3200 0.7050 0.6950 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8950 0.3500 1.6500 ;
        RECT 0.2500 1.6500 0.7450 1.7500 ;
        RECT 0.2500 0.7950 0.4500 0.8950 ;
        RECT 0.5750 1.7500 0.7450 1.9600 ;
        RECT 0.3500 0.5000 0.4500 0.7950 ;
    END
    ANTENNADIFFAREA 0.20125 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0550 1.8550 0.2250 2.0800 ;
    END
  END VDD
END NOR2_X1B_A12TH

MACRO NOR2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6700 ;
        RECT 0.6150 0.3200 0.7050 0.8600 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8950 0.3500 1.6500 ;
        RECT 0.2500 1.6500 0.7450 1.7500 ;
        RECT 0.2500 0.7950 0.4500 0.8950 ;
        RECT 0.5750 1.7500 0.7450 1.9600 ;
        RECT 0.3500 0.4250 0.4500 0.7950 ;
    END
    ANTENNADIFFAREA 0.23425 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0550 1.8550 0.2250 2.0800 ;
    END
  END VDD
END NOR2_X1M_A12TH

MACRO NOR2_X1P4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7650 ;
        RECT 0.6100 0.3200 0.7100 0.5500 ;
        RECT 1.1300 0.3200 1.2300 0.5500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.2500 1.1500 1.3500 ;
        RECT 1.0500 1.0500 1.1500 1.2500 ;
        RECT 0.1950 0.8900 0.2950 1.2500 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0500 0.8700 1.1500 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.4500 1.3500 1.5500 ;
        RECT 0.6100 1.5500 0.7100 1.8900 ;
        RECT 1.2500 0.7500 1.3500 1.4500 ;
        RECT 0.3150 0.6500 1.3500 0.7500 ;
        RECT 0.3150 0.4400 0.4850 0.6500 ;
        RECT 0.8350 0.4400 1.0050 0.6500 ;
    END
    ANTENNADIFFAREA 0.291 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1300 1.6450 1.2300 2.0800 ;
        RECT 0.0900 1.5900 0.1900 2.0800 ;
    END
  END VDD
END NOR2_X1P4A_A12TH

MACRO NOR2_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5400 ;
        RECT 0.5950 0.3200 0.6950 0.5400 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 1.0300 0.7950 1.1500 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.2500 1.0200 1.3500 ;
        RECT 0.9200 1.0200 1.0200 1.2500 ;
        RECT 0.2350 1.0100 0.3350 1.2500 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0550 1.4500 0.6600 1.5500 ;
        RECT 0.5700 1.5500 0.6600 1.9850 ;
        RECT 0.0550 0.7600 0.1450 1.4500 ;
        RECT 0.0550 0.6700 0.4350 0.7600 ;
        RECT 0.3350 0.4700 0.4350 0.6700 ;
    END
    ANTENNADIFFAREA 0.199 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.0750 1.7550 0.1750 2.0800 ;
        RECT 1.0250 1.7550 1.1250 2.0800 ;
    END
  END VDD
END NOR2_X1P4B_A12TH

MACRO NOR2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0850 0.3200 0.1750 0.8000 ;
        RECT 0.6050 0.3200 0.6950 0.8000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.0850 1.7300 0.1750 2.0800 ;
        RECT 1.0300 1.7300 1.1200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4500 0.6700 1.5500 ;
        RECT 0.5800 1.5500 0.6700 1.9800 ;
        RECT 0.0500 0.9800 0.1500 1.4500 ;
        RECT 0.0500 0.8900 0.4350 0.9800 ;
        RECT 0.3450 0.4950 0.4350 0.8900 ;
    END
    ANTENNADIFFAREA 0.235 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 1.1050 1.3500 ;
        RECT 0.9150 1.3500 1.1050 1.3750 ;
        RECT 0.2400 1.1300 0.3400 1.2500 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5250 1.0500 0.9450 1.1500 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END A
END NOR2_X1P4M_A12TH

MACRO NOR2_X2A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7400 ;
        RECT 0.5800 0.3200 0.7500 0.6300 ;
        RECT 1.1000 0.3200 1.2700 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.4500 1.1500 1.5500 ;
        RECT 0.1950 0.9800 0.2950 1.4500 ;
        RECT 1.0500 0.9800 1.1500 1.4500 ;
    END
    ANTENNAGATEAREA 0.1776 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.1776 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5800 1.6500 1.3500 1.7500 ;
        RECT 0.5800 1.7500 0.7500 1.9700 ;
        RECT 1.2500 0.8400 1.3500 1.6500 ;
        RECT 0.3550 0.7400 1.3500 0.8400 ;
        RECT 0.8750 0.4200 0.9750 0.7400 ;
        RECT 0.3550 0.4100 0.4550 0.7400 ;
    END
    ANTENNADIFFAREA 0.41 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1000 1.8600 1.2700 2.0800 ;
        RECT 0.0950 1.7700 0.1950 2.0800 ;
    END
  END VDD
END NOR2_X2A_A12TH

MACRO NOR2_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5800 ;
        RECT 0.5950 0.3200 0.6950 0.6100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 1.0300 0.7950 1.1500 ;
    END
    ANTENNAGATEAREA 0.1344 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.2500 1.0200 1.3500 ;
        RECT 0.9200 1.0200 1.0200 1.2500 ;
        RECT 0.2350 1.0100 0.3350 1.2500 ;
    END
    ANTENNAGATEAREA 0.1344 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0550 1.4500 0.6600 1.5500 ;
        RECT 0.5700 1.5500 0.6600 1.8900 ;
        RECT 0.0550 0.7600 0.1450 1.4500 ;
        RECT 0.0550 0.6700 0.4350 0.7600 ;
        RECT 0.3350 0.4100 0.4350 0.6700 ;
    END
    ANTENNADIFFAREA 0.266 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.0750 1.7550 0.1750 2.0800 ;
        RECT 1.0250 1.7550 1.1250 2.0800 ;
    END
  END VDD
END NOR2_X2B_A12TH

MACRO NOR2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5800 ;
        RECT 0.6000 0.3200 0.6900 0.6100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 1.0300 0.7950 1.1500 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.2500 1.0200 1.3500 ;
        RECT 0.9200 1.0200 1.0200 1.2500 ;
        RECT 0.2350 1.0100 0.3350 1.2500 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0550 1.4500 0.6600 1.5500 ;
        RECT 0.5700 1.5500 0.6600 1.8900 ;
        RECT 0.0550 0.7600 0.1450 1.4500 ;
        RECT 0.0550 0.6700 0.4700 0.7600 ;
        RECT 0.3000 0.4100 0.4700 0.6700 ;
    END
    ANTENNADIFFAREA 0.332 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.0800 1.7550 0.1700 2.0800 ;
        RECT 1.0300 1.7550 1.1200 2.0800 ;
    END
  END VDD
END NOR2_X2M_A12TH

MACRO NOR2_X3A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.6150 ;
        RECT 0.6050 0.3200 0.7750 0.5100 ;
        RECT 1.1250 0.3200 1.2950 0.5100 ;
        RECT 1.6450 0.3200 1.8150 0.5100 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 1.4000 1.1500 ;
    END
    ANTENNAGATEAREA 0.2664 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 0.8500 1.6150 0.9500 ;
        RECT 1.5150 0.9500 1.6150 1.1000 ;
    END
    ANTENNAGATEAREA 0.2664 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 1.4500 1.9500 1.5500 ;
        RECT 0.6400 1.5500 0.7400 1.8800 ;
        RECT 1.6800 1.5500 1.7800 1.8800 ;
        RECT 1.8500 0.7500 1.9500 1.4500 ;
        RECT 0.3450 0.6500 1.9500 0.7500 ;
        RECT 0.3450 0.4400 0.5150 0.6500 ;
        RECT 0.8650 0.4400 1.0350 0.6500 ;
        RECT 1.3850 0.4400 1.5550 0.6500 ;
    END
    ANTENNADIFFAREA 0.7151 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1200 1.7550 0.2200 2.0800 ;
        RECT 1.1600 1.7550 1.2600 2.0800 ;
    END
  END VDD
END NOR2_X3A_A12TH

MACRO NOR2_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3900 0.3200 0.4800 0.5600 ;
        RECT 0.9800 0.3200 1.0700 0.5600 ;
        RECT 1.5800 0.3200 1.6700 0.6450 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.5900 1.7550 0.6800 2.0800 ;
        RECT 1.5900 1.7550 1.6800 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.2500 1.5650 1.3500 ;
        RECT 0.7500 1.2150 0.8500 1.2500 ;
        RECT 1.4650 1.2000 1.5650 1.2500 ;
        RECT 0.4600 1.1150 0.8500 1.2150 ;
        RECT 1.4650 1.1000 1.6650 1.2000 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.6500 1.4500 0.7500 ;
        RECT 0.0450 0.7500 0.1350 1.5100 ;
        RECT 0.6100 0.5400 0.7800 0.6500 ;
        RECT 1.2800 0.5400 1.4500 0.6500 ;
        RECT 0.0450 1.5100 1.1900 1.6000 ;
        RECT 0.0450 1.6000 0.1700 1.9500 ;
        RECT 1.1000 1.6000 1.1900 1.9500 ;
    END
    ANTENNADIFFAREA 0.4536 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8450 1.2250 0.9500 ;
        RECT 0.2350 0.9500 0.3250 1.0500 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END A
END NOR2_X3B_A12TH

MACRO NOR2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.3900 0.3200 0.4800 0.5600 ;
        RECT 0.9800 0.3200 1.0700 0.5600 ;
        RECT 1.5800 0.3200 1.6700 0.6450 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.5900 1.7550 0.6800 2.0800 ;
        RECT 1.5900 1.7550 1.6800 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.2500 1.5650 1.3500 ;
        RECT 0.7500 1.2150 0.8500 1.2500 ;
        RECT 1.4650 1.2000 1.5650 1.2500 ;
        RECT 0.4600 1.1150 0.8500 1.2150 ;
        RECT 1.4650 1.1000 1.6650 1.2000 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.6500 1.4500 0.7500 ;
        RECT 0.0450 0.7500 0.1350 1.5100 ;
        RECT 0.6100 0.4100 0.7800 0.6500 ;
        RECT 1.2800 0.4100 1.4500 0.6500 ;
        RECT 0.0450 1.5100 1.1900 1.6000 ;
        RECT 0.0450 1.6000 0.1700 1.9500 ;
        RECT 1.1000 1.6000 1.1900 1.9500 ;
    END
    ANTENNADIFFAREA 0.5536 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8450 1.2250 0.9500 ;
        RECT 0.2350 0.9500 0.3250 1.0500 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END A
END NOR2_X3M_A12TH

MACRO NOR2_X4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 1.0350 1.7700 1.1350 2.0800 ;
        RECT 2.0250 1.7700 2.1250 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.4650 0.3200 0.5650 0.6400 ;
        RECT 0.9850 0.3200 1.0850 0.5600 ;
        RECT 1.5050 0.3200 1.6050 0.5600 ;
        RECT 2.0250 0.3200 2.1250 0.5400 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1450 0.8500 1.9500 0.9500 ;
        RECT 1.1450 0.9500 1.2450 1.0500 ;
        RECT 1.8500 0.9500 1.9500 1.2350 ;
        RECT 0.8550 1.0500 1.2450 1.1500 ;
        RECT 0.8550 0.9500 0.9550 1.0500 ;
        RECT 0.1800 0.8500 0.9550 0.9500 ;
        RECT 0.1800 0.9500 0.2800 1.2200 ;
    END
    ANTENNAGATEAREA 0.3552 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6750 1.2500 1.4450 1.3500 ;
        RECT 0.6750 1.1900 0.7650 1.2500 ;
        RECT 1.3550 1.1850 1.4450 1.2500 ;
        RECT 0.3950 1.0900 0.7650 1.1900 ;
        RECT 1.3550 1.0850 1.7400 1.1850 ;
    END
    ANTENNAGATEAREA 0.3552 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.7500 2.1500 1.4500 ;
        RECT 0.5350 1.4500 2.1500 1.5500 ;
        RECT 0.6900 0.6500 2.1500 0.7500 ;
        RECT 0.5350 1.5500 0.6350 1.8700 ;
        RECT 1.5050 1.5500 1.6050 1.8800 ;
        RECT 0.6900 0.4550 0.8600 0.6500 ;
        RECT 1.2100 0.4550 1.3800 0.6500 ;
        RECT 1.7300 0.4550 1.9000 0.6500 ;
    END
    ANTENNADIFFAREA 0.82 ;
  END Y
END NOR2_X4A_A12TH

MACRO NOR2_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 1.0450 1.7700 1.1450 2.0800 ;
        RECT 2.0250 1.7700 2.1250 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.7250 0.3200 0.8250 0.5250 ;
        RECT 1.2450 0.3200 1.3450 0.5250 ;
        RECT 1.7650 0.3200 1.8650 0.5250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1250 0.8500 1.9550 0.9500 ;
        RECT 1.8550 0.9500 1.9550 1.1900 ;
    END
    ANTENNAGATEAREA 0.2688 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4050 1.0500 1.7450 1.1500 ;
    END
    ANTENNAGATEAREA 0.2688 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.7500 2.1500 1.4500 ;
        RECT 0.5350 1.4500 2.1500 1.5500 ;
        RECT 0.9500 0.6500 2.1500 0.7500 ;
        RECT 0.5350 1.5500 0.6350 1.8800 ;
        RECT 1.5050 1.5500 1.6050 1.8800 ;
        RECT 1.4700 0.4250 1.6400 0.6500 ;
        RECT 0.9500 0.4100 1.1200 0.6500 ;
    END
    ANTENNADIFFAREA 0.532 ;
  END Y
END NOR2_X4B_A12TH

MACRO NOR2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.4650 0.3200 0.5650 0.6500 ;
        RECT 0.9850 0.3200 1.0850 0.4450 ;
        RECT 1.5050 0.3200 1.6050 0.4450 ;
        RECT 2.0250 0.3200 2.1250 0.4450 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1800 0.8500 1.9550 0.9500 ;
        RECT 0.1800 0.9500 0.2800 1.1900 ;
        RECT 1.8550 0.9500 1.9550 1.1900 ;
    END
    ANTENNAGATEAREA 0.3084 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4050 1.0500 1.7450 1.1500 ;
    END
    ANTENNAGATEAREA 0.3084 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.7500 2.1500 1.4500 ;
        RECT 0.5350 1.4500 2.1500 1.5500 ;
        RECT 0.6900 0.6500 2.1500 0.7500 ;
        RECT 0.5350 1.5500 0.6350 1.8800 ;
        RECT 1.5050 1.5500 1.6050 1.8800 ;
        RECT 0.6900 0.4250 0.8600 0.6500 ;
        RECT 1.2100 0.4250 1.3800 0.6500 ;
        RECT 1.7300 0.4250 1.9000 0.6500 ;
    END
    ANTENNADIFFAREA 0.664 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 1.0450 1.7700 1.1450 2.0800 ;
        RECT 2.0250 1.7700 2.1250 2.0800 ;
    END
  END VDD
END NOR2_X4M_A12TH

MACRO NOR2_X6A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0850 0.3200 0.1750 0.5800 ;
        RECT 0.6000 0.3200 0.7000 0.5600 ;
        RECT 1.1200 0.3200 1.2200 0.5600 ;
        RECT 1.6400 0.3200 1.7400 0.5600 ;
        RECT 2.1650 0.3200 2.2650 0.5600 ;
        RECT 2.6850 0.3200 2.7850 0.5600 ;
        RECT 3.2050 0.3200 3.3050 0.5600 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1800 1.0500 3.1550 1.1500 ;
    END
    ANTENNAGATEAREA 0.5328 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 0.8500 2.9000 0.9500 ;
    END
    ANTENNAGATEAREA 0.5328 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6000 1.4500 3.3500 1.5500 ;
        RECT 0.6000 1.5500 0.7000 1.8850 ;
        RECT 1.6400 1.5500 1.7400 1.8850 ;
        RECT 2.6850 1.5500 2.7850 1.8850 ;
        RECT 3.2500 0.7500 3.3500 1.4500 ;
        RECT 0.3050 0.6500 3.3500 0.7500 ;
        RECT 0.3050 0.4400 0.4750 0.6500 ;
        RECT 0.8250 0.4400 0.9950 0.6500 ;
        RECT 1.3450 0.4400 1.5150 0.6500 ;
        RECT 1.8700 0.4400 2.0400 0.6500 ;
        RECT 2.3900 0.4400 2.5600 0.6500 ;
        RECT 2.9100 0.4400 3.0800 0.6500 ;
    END
    ANTENNADIFFAREA 1.23455 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0800 1.7650 0.1800 2.0800 ;
        RECT 1.1200 1.7650 1.2200 2.0800 ;
        RECT 2.1650 1.7650 2.2650 2.0800 ;
        RECT 3.2050 1.7650 3.3050 2.0800 ;
    END
  END VDD
END NOR2_X6A_A12TH

MACRO NOR2_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 1.2500 0.3200 1.3400 0.6000 ;
        RECT 1.7700 0.3200 1.8600 0.6000 ;
        RECT 2.2900 0.3200 2.3800 0.6000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.2500 2.4250 1.3500 ;
        RECT 2.3350 1.1800 2.4250 1.2500 ;
        RECT 1.3650 1.0700 1.7350 1.2500 ;
        RECT 0.4100 1.0500 0.5550 1.2500 ;
        RECT 2.3350 1.0900 2.7250 1.1800 ;
    END
    ANTENNAGATEAREA 0.4032 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.2550 1.1500 ;
        RECT 1.1600 0.9600 1.2550 1.0500 ;
        RECT 1.1600 0.8700 2.9750 0.9600 ;
        RECT 1.8450 0.9600 1.9350 1.0700 ;
        RECT 1.8450 1.0700 2.2250 1.1600 ;
    END
    ANTENNAGATEAREA 0.4032 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.4500 2.5600 1.5500 ;
        RECT 0.5400 1.5500 0.6300 1.8800 ;
        RECT 1.5100 1.5500 1.6000 1.8700 ;
        RECT 2.4700 1.5500 2.5600 1.8700 ;
        RECT 0.2300 0.7800 0.3200 1.4500 ;
        RECT 0.2300 0.6900 2.1200 0.7800 ;
        RECT 1.5100 0.4100 1.6000 0.6900 ;
        RECT 2.0300 0.4100 2.1200 0.6900 ;
    END
    ANTENNADIFFAREA 0.798 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0800 1.7450 0.1700 2.0800 ;
        RECT 1.0250 1.7450 1.1150 2.0800 ;
        RECT 1.9950 1.7450 2.0850 2.0800 ;
        RECT 2.9300 1.7450 3.0200 2.0800 ;
    END
  END VDD
END NOR2_X6B_A12TH

MACRO NOR2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.9900 0.3200 1.0800 0.6000 ;
        RECT 1.5100 0.3200 1.6000 0.6000 ;
        RECT 2.0300 0.3200 2.1200 0.6000 ;
        RECT 2.5500 0.3200 2.6400 0.6000 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.2550 1.1500 ;
        RECT 1.1600 0.9600 1.2550 1.0500 ;
        RECT 1.1600 0.8700 2.9800 0.9600 ;
        RECT 1.8450 0.9600 1.9350 1.0700 ;
        RECT 1.8450 1.0700 2.2250 1.1600 ;
    END
    ANTENNAGATEAREA 0.4626 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.4500 2.5600 1.5500 ;
        RECT 0.5400 1.5500 0.6300 1.8800 ;
        RECT 1.5100 1.5500 1.6000 1.8700 ;
        RECT 2.4700 1.5500 2.5600 1.8700 ;
        RECT 0.2300 0.7800 0.3200 1.4500 ;
        RECT 0.2300 0.6900 2.3800 0.7800 ;
        RECT 1.2500 0.4100 1.3400 0.6900 ;
        RECT 1.7700 0.4100 1.8600 0.6900 ;
        RECT 2.2900 0.4100 2.3800 0.6900 ;
    END
    ANTENNADIFFAREA 0.996 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.2500 2.4250 1.3500 ;
        RECT 2.3350 1.1800 2.4250 1.2500 ;
        RECT 1.3650 1.0700 1.7350 1.2500 ;
        RECT 0.4100 1.0500 0.5550 1.2500 ;
        RECT 2.3350 1.0900 2.7250 1.1800 ;
    END
    ANTENNAGATEAREA 0.4626 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0800 1.7450 0.1700 2.0800 ;
        RECT 1.0250 1.7450 1.1150 2.0800 ;
        RECT 1.9950 1.7450 2.0850 2.0800 ;
        RECT 2.9300 1.7450 3.0200 2.0800 ;
    END
  END VDD
END NOR2_X6M_A12TH

MACRO NOR2_X8A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1900 0.3200 0.2900 0.6300 ;
        RECT 0.6750 0.3200 0.8450 0.5250 ;
        RECT 1.1950 0.3200 1.3650 0.5250 ;
        RECT 1.7200 0.3200 1.8900 0.5250 ;
        RECT 2.2400 0.3200 2.4100 0.5250 ;
        RECT 2.7600 0.3200 2.9300 0.5250 ;
        RECT 3.2800 0.3200 3.4500 0.5250 ;
        RECT 3.8000 0.3200 3.9700 0.5250 ;
        RECT 4.3200 0.3200 4.4900 0.5250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 4.3000 1.1500 ;
        RECT 4.2000 0.9450 4.3000 1.0500 ;
    END
    ANTENNAGATEAREA 0.7104 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5700 0.8500 4.0400 0.9500 ;
    END
    ANTENNAGATEAREA 0.7104 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7100 1.4350 4.5500 1.5650 ;
        RECT 0.7100 1.5650 0.8100 1.8650 ;
        RECT 1.7500 1.5650 1.8500 1.8650 ;
        RECT 2.7950 1.5650 2.8950 1.8650 ;
        RECT 3.8350 1.5650 3.9350 1.8650 ;
        RECT 4.4200 0.7500 4.5500 1.4350 ;
        RECT 0.4150 0.6200 4.5500 0.7500 ;
        RECT 0.4150 0.4200 0.5850 0.6200 ;
        RECT 0.9350 0.4200 1.1050 0.6200 ;
        RECT 1.4550 0.4200 1.6250 0.6200 ;
        RECT 1.9800 0.4200 2.1500 0.6200 ;
        RECT 2.5000 0.4200 2.6700 0.6200 ;
        RECT 3.0200 0.4200 3.1900 0.6200 ;
        RECT 3.5400 0.4200 3.7100 0.6200 ;
        RECT 4.0600 0.4200 4.2300 0.6200 ;
    END
    ANTENNADIFFAREA 1.64455 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1900 1.7700 0.2900 2.0800 ;
        RECT 1.2300 1.7700 1.3300 2.0800 ;
        RECT 2.2750 1.7700 2.3750 2.0800 ;
        RECT 3.3150 1.7700 3.4150 2.0800 ;
        RECT 4.3550 1.7700 4.4550 2.0800 ;
    END
  END VDD
END NOR2_X8A_A12TH

MACRO NOR2_X8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1900 0.3200 0.2900 0.5700 ;
        RECT 0.6750 0.3200 0.8450 0.5250 ;
        RECT 1.1950 0.3200 1.3650 0.5250 ;
        RECT 1.7200 0.3200 1.8900 0.5250 ;
        RECT 2.2400 0.3200 2.4100 0.5250 ;
        RECT 2.7600 0.3200 2.9300 0.5250 ;
        RECT 3.2800 0.3200 3.4500 0.5250 ;
        RECT 3.8000 0.3200 3.9700 0.5250 ;
        RECT 4.3200 0.3200 4.4900 0.5250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 4.3000 1.1500 ;
        RECT 4.2000 0.9450 4.3000 1.0500 ;
    END
    ANTENNAGATEAREA 0.5376 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5700 0.8500 4.0400 0.9500 ;
    END
    ANTENNAGATEAREA 0.5376 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7100 1.4350 4.5500 1.5650 ;
        RECT 0.7100 1.5650 0.8100 1.8650 ;
        RECT 1.7500 1.5650 1.8500 1.8650 ;
        RECT 2.7950 1.5650 2.8950 1.8650 ;
        RECT 3.8350 1.5650 3.9350 1.8650 ;
        RECT 4.4200 0.7500 4.5500 1.4350 ;
        RECT 0.4150 0.6200 4.5500 0.7500 ;
        RECT 0.4150 0.4200 0.5850 0.6200 ;
        RECT 0.9350 0.4200 1.1050 0.6200 ;
        RECT 1.4550 0.4200 1.6250 0.6200 ;
        RECT 1.9800 0.4200 2.1500 0.6200 ;
        RECT 2.5000 0.4200 2.6700 0.6200 ;
        RECT 3.0200 0.4200 3.1900 0.6200 ;
        RECT 3.5400 0.4200 3.7100 0.6200 ;
        RECT 4.0600 0.4200 4.2300 0.6200 ;
    END
    ANTENNADIFFAREA 1.06855 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1900 1.7700 0.2900 2.0800 ;
        RECT 1.2300 1.7700 1.3300 2.0800 ;
        RECT 2.2750 1.7700 2.3750 2.0800 ;
        RECT 3.3150 1.7700 3.4150 2.0800 ;
        RECT 4.3550 1.7700 4.4550 2.0800 ;
    END
  END VDD
END NOR2_X8B_A12TH

MACRO NOR2_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1900 0.3200 0.2900 0.8000 ;
        RECT 0.6750 0.3200 0.8450 0.4950 ;
        RECT 1.1950 0.3200 1.3650 0.4950 ;
        RECT 1.7200 0.3200 1.8900 0.4950 ;
        RECT 2.2400 0.3200 2.4100 0.4950 ;
        RECT 2.7600 0.3200 2.9300 0.4950 ;
        RECT 3.2800 0.3200 3.4500 0.4950 ;
        RECT 3.8000 0.3200 3.9700 0.4950 ;
        RECT 4.3200 0.3200 4.4900 0.4950 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 4.3000 1.1500 ;
        RECT 4.2000 0.9450 4.3000 1.0500 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5700 0.8500 4.0400 0.9500 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7100 1.4350 4.5500 1.5650 ;
        RECT 0.7100 1.5650 0.8100 1.8650 ;
        RECT 1.7500 1.5650 1.8500 1.8650 ;
        RECT 2.7950 1.5650 2.8950 1.8650 ;
        RECT 3.8350 1.5650 3.9350 1.8650 ;
        RECT 4.4200 0.7500 4.5500 1.4350 ;
        RECT 0.4150 0.6200 4.5500 0.7500 ;
        RECT 0.4150 0.4200 0.5850 0.6200 ;
        RECT 0.9350 0.4200 1.1050 0.6200 ;
        RECT 1.4550 0.4200 1.6250 0.6200 ;
        RECT 1.9800 0.4200 2.1500 0.6200 ;
        RECT 2.5000 0.4200 2.6700 0.6200 ;
        RECT 3.0200 0.4200 3.1900 0.6200 ;
        RECT 3.5400 0.4200 3.7100 0.6200 ;
        RECT 4.0600 0.4200 4.2300 0.6200 ;
    END
    ANTENNADIFFAREA 1.33255 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1900 1.7700 0.2900 2.0800 ;
        RECT 1.2300 1.7700 1.3300 2.0800 ;
        RECT 2.2750 1.7700 2.3750 2.0800 ;
        RECT 3.3150 1.7700 3.4150 2.0800 ;
        RECT 4.3550 1.7700 4.4550 2.0800 ;
    END
  END VDD
END NOR2_X8M_A12TH

MACRO NOR3_X0P5A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6950 ;
        RECT 0.8700 0.3200 0.9700 0.6950 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9950 0.3500 1.4150 ;
    END
    ANTENNAGATEAREA 0.0405 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1000 0.5500 1.3900 ;
        RECT 0.4500 1.0000 0.7000 1.1000 ;
    END
    ANTENNAGATEAREA 0.0405 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8850 0.1500 1.5100 ;
        RECT 0.0500 1.5100 0.1850 1.9000 ;
        RECT 0.0500 0.7850 0.7100 0.8850 ;
        RECT 0.0500 0.5050 0.1700 0.7850 ;
        RECT 0.6100 0.5000 0.7100 0.7850 ;
    END
    ANTENNADIFFAREA 0.162125 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.8700 1.5000 0.9700 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8900 0.9600 1.3050 ;
    END
    ANTENNAGATEAREA 0.0405 ;
  END C
END NOR3_X0P5A_A12TH

MACRO NOR3_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7100 ;
        RECT 0.8700 0.3200 0.9700 0.7100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.3900 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1000 0.5500 1.3900 ;
        RECT 0.4500 1.0000 0.7000 1.1000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9000 0.1500 1.4700 ;
        RECT 0.0500 1.4700 0.1900 1.8600 ;
        RECT 0.0500 0.8000 0.7100 0.9000 ;
        RECT 0.0950 0.5200 0.1850 0.8000 ;
        RECT 0.6100 0.5150 0.7100 0.8000 ;
    END
    ANTENNADIFFAREA 0.1525 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.8700 1.4950 0.9700 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8900 0.9600 1.3050 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END C
END NOR3_X0P5M_A12TH

MACRO NOR3_X0P7A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7100 ;
        RECT 0.8550 0.3200 0.9550 0.7350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.5400 0.2200 1.8300 ;
        RECT 0.0500 0.9000 0.1500 1.5400 ;
        RECT 0.0500 0.8000 0.6950 0.9000 ;
        RECT 0.0500 0.6450 0.1700 0.8000 ;
        RECT 0.5950 0.6450 0.6950 0.8000 ;
    END
    ANTENNADIFFAREA 0.256725 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0573 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 0.9100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0573 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.0500 1.1250 1.1500 ;
    END
    ANTENNAGATEAREA 0.0573 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.8550 1.6800 0.9550 2.0800 ;
    END
  END VDD
END NOR3_X0P7A_A12TH

MACRO NOR3_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7100 ;
        RECT 0.8700 0.3200 0.9700 0.7100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.8700 1.5450 0.9700 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8900 0.9600 1.3050 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1000 0.5500 1.3900 ;
        RECT 0.4500 1.0000 0.7000 1.1000 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9000 0.1500 1.5100 ;
        RECT 0.0500 1.5100 0.1900 1.9000 ;
        RECT 0.0500 0.8000 0.7100 0.9000 ;
        RECT 0.0950 0.5200 0.1850 0.8000 ;
        RECT 0.6100 0.5150 0.7100 0.8000 ;
    END
    ANTENNADIFFAREA 0.1785 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END A
END NOR3_X0P7M_A12TH

MACRO NOR3_X1A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4600 0.3200 0.5600 0.7100 ;
        RECT 0.9800 0.3200 1.0800 0.7650 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9000 0.1500 1.5400 ;
        RECT 0.0500 1.5400 0.2250 1.9700 ;
        RECT 0.0500 0.8000 0.8200 0.9000 ;
        RECT 0.0500 0.4450 0.1700 0.8000 ;
        RECT 0.7200 0.4400 0.8200 0.8000 ;
    END
    ANTENNADIFFAREA 0.44575 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4300 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9900 0.7550 1.4250 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.9450 1.1500 1.3650 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9800 1.7700 1.0800 2.0800 ;
    END
  END VDD
END NOR3_X1A_A12TH

MACRO NOR3_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7050 ;
        RECT 0.8700 0.3200 0.9700 0.7050 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1000 0.5500 1.3900 ;
        RECT 0.4500 1.0000 0.7000 1.1000 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8900 0.9600 1.3050 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9000 0.1500 1.4700 ;
        RECT 0.0500 1.4700 0.1900 1.8600 ;
        RECT 0.0500 0.8000 0.7100 0.9000 ;
        RECT 0.0950 0.5200 0.1850 0.8000 ;
        RECT 0.6100 0.5150 0.7100 0.8000 ;
    END
    ANTENNADIFFAREA 0.253 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.8700 1.7900 0.9700 2.0800 ;
    END
  END VDD
END NOR3_X1M_A12TH

MACRO NAND4_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 2.2150 0.3200 2.3850 0.5300 ;
        RECT 3.2550 0.3200 3.4250 0.5250 ;
        RECT 4.2100 0.3200 4.3100 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4050 1.0450 1.7350 1.1550 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1850 1.4500 3.1300 1.5500 ;
        RECT 1.1850 1.5500 1.2850 1.9000 ;
        RECT 1.7350 1.5500 1.8350 1.9000 ;
        RECT 2.5100 1.5500 2.6100 1.9000 ;
        RECT 3.0300 1.5500 3.1300 1.9000 ;
        RECT 2.0850 0.9500 2.1850 1.4500 ;
        RECT 0.5550 0.8500 2.1850 0.9500 ;
        RECT 0.5550 0.7100 0.6550 0.8500 ;
        RECT 1.4750 0.7100 1.5750 0.8500 ;
    END
    ANTENNADIFFAREA 0.93215 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2950 1.2500 3.5000 1.3500 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6200 1.0500 3.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8350 1.2500 1.9750 1.3500 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 0.8950 1.7700 0.9950 2.0800 ;
        RECT 1.4750 1.7700 1.5750 2.0800 ;
        RECT 1.9950 1.7700 2.0950 2.0800 ;
        RECT 2.2500 1.7700 2.3500 2.0800 ;
        RECT 2.7700 1.7700 2.8700 2.0800 ;
        RECT 3.2900 1.7700 3.3900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.9400 0.6650 3.8850 0.7550 ;
      RECT 3.7150 0.4250 3.8850 0.6650 ;
      RECT 0.0800 0.4800 2.0300 0.5700 ;
      RECT 1.9400 0.5700 2.0300 0.6650 ;
      RECT 0.0800 0.5700 0.1700 0.9100 ;
      RECT 2.7350 0.4250 2.9050 0.6650 ;
  END
END NAND4_X4M_A12TH

MACRO NOR2B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4200 0.3200 0.5200 0.6000 ;
        RECT 0.9850 0.3200 1.1550 0.5050 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7500 0.3500 1.1700 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 0.8050 0.7500 1.2150 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7000 1.1500 1.6850 ;
        RECT 0.9750 1.6850 1.1500 1.9800 ;
        RECT 0.7500 0.6100 1.1500 0.7000 ;
        RECT 0.7500 0.4100 0.8500 0.6100 ;
    END
    ANTENNADIFFAREA 0.120325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3750 1.6900 0.5450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.5000 0.9500 1.5900 ;
      RECT 0.8600 1.0000 0.9500 1.5000 ;
      RECT 0.0550 0.4500 0.2500 0.5400 ;
      RECT 0.0550 1.5900 0.1850 1.7400 ;
      RECT 0.0550 0.5400 0.1450 1.5000 ;
  END
END NOR2B_X0P5M_A12TH

MACRO NOR2B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4200 0.3200 0.5200 0.6250 ;
        RECT 0.9850 0.3200 1.1550 0.4950 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 0.8400 0.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7500 0.3500 1.1800 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.6900 1.1500 1.6600 ;
        RECT 0.9750 1.6600 1.1500 1.9800 ;
        RECT 0.7500 0.5900 1.1500 0.6900 ;
        RECT 0.7500 0.4200 0.8500 0.5900 ;
    END
    ANTENNADIFFAREA 0.171175 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4400 1.7650 0.5500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.4600 0.9500 1.5500 ;
      RECT 0.8600 0.8950 0.9500 1.4600 ;
      RECT 0.0550 0.4700 0.2500 0.5700 ;
      RECT 0.0550 1.5500 0.1850 1.7400 ;
      RECT 0.0550 0.5700 0.1450 1.4600 ;
  END
END NOR2B_X0P7M_A12TH

MACRO NOR2B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4350 0.3200 0.5350 0.8200 ;
        RECT 0.9250 0.3200 1.0950 0.7200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.5400 ;
        RECT 0.9800 1.5400 1.1500 1.6400 ;
        RECT 0.6950 0.8500 1.1500 0.9500 ;
        RECT 0.9800 1.6400 1.0800 1.9600 ;
        RECT 0.6950 0.4200 0.7950 0.8500 ;
    END
    ANTENNADIFFAREA 0.2752 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.1500 0.3500 1.5950 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9300 0.5500 1.3550 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4000 1.8950 0.5700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.7050 0.8750 1.7950 ;
      RECT 0.7850 1.0500 0.8750 1.7050 ;
      RECT 0.0500 0.6600 0.2500 0.7500 ;
      RECT 0.0500 0.7500 0.1400 1.7050 ;
  END
END NOR2B_X1M_A12TH

MACRO NOR2B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3600 0.3200 0.4700 0.5200 ;
        RECT 0.8800 0.3200 0.9900 0.5300 ;
        RECT 1.4000 0.3200 1.5100 0.5300 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7650 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0333 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7500 1.5500 1.4500 ;
        RECT 0.8850 1.4500 1.5500 1.5500 ;
        RECT 0.6250 0.6500 1.5500 0.7500 ;
        RECT 0.8850 1.5500 0.9850 1.9000 ;
        RECT 0.6250 0.4250 0.7250 0.6500 ;
        RECT 1.1450 0.4250 1.2450 0.6500 ;
    END
    ANTENNADIFFAREA 0.235 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.4050 1.6700 1.5050 2.0800 ;
        RECT 0.4050 1.6350 0.5050 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 0.8500 1.3350 0.9500 ;
        RECT 1.2350 0.9500 1.3350 1.0600 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.7100 1.0950 1.1250 1.1850 ;
      RECT 0.0550 0.4100 0.2500 0.5000 ;
      RECT 0.0550 1.3900 0.1750 1.6150 ;
      RECT 0.0550 0.5000 0.1450 1.3000 ;
      RECT 0.0550 1.3000 0.8000 1.3900 ;
      RECT 0.7100 1.1850 0.8000 1.3000 ;
  END
END NOR2B_X1P4M_A12TH

MACRO NOR2B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3300 0.3200 0.5000 0.6150 ;
        RECT 0.8800 0.3200 0.9900 0.4550 ;
        RECT 1.4000 0.3200 1.5100 0.4550 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7650 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7500 1.5500 1.4500 ;
        RECT 0.8850 1.4500 1.5500 1.5500 ;
        RECT 0.6250 0.6500 1.5500 0.7500 ;
        RECT 0.8850 1.5500 0.9850 1.8900 ;
        RECT 0.6250 0.4350 0.7250 0.6500 ;
        RECT 1.1450 0.4300 1.2450 0.6500 ;
    END
    ANTENNADIFFAREA 0.332 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4750 0.8500 1.3350 0.9500 ;
        RECT 1.2350 0.9500 1.3350 1.0600 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3550 1.7700 0.4550 2.0800 ;
        RECT 1.4050 1.7700 1.5050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.1250 1.1500 ;
      RECT 0.0550 1.5000 0.7900 1.5900 ;
      RECT 0.7000 1.1500 0.7900 1.5000 ;
      RECT 0.0550 1.5900 0.1850 1.9700 ;
      RECT 0.0550 0.5550 0.1450 1.5000 ;
      RECT 0.0550 0.4650 0.2400 0.5550 ;
  END
END NOR2B_X2M_A12TH

MACRO NOR2B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.5050 0.3200 0.6050 0.5600 ;
        RECT 1.0300 0.3200 1.1300 0.5600 ;
        RECT 1.5500 0.3200 1.6500 0.5950 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 0.8500 1.5300 0.9600 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.7950 1.7500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0648 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7500 0.1500 1.4500 ;
        RECT 0.0500 1.4500 1.1300 1.5500 ;
        RECT 0.0500 0.6500 1.3900 0.7500 ;
        RECT 0.0500 1.5500 0.1700 1.9150 ;
        RECT 1.0300 1.5500 1.1300 1.9200 ;
        RECT 0.7700 0.5200 0.8700 0.6500 ;
        RECT 1.2900 0.5000 1.3900 0.6500 ;
    END
    ANTENNADIFFAREA 0.556425 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.5700 1.7700 0.6700 2.0800 ;
        RECT 1.5500 1.6800 1.6500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.8300 1.5800 1.9450 1.9550 ;
      RECT 1.2300 1.4900 1.9450 1.5800 ;
      RECT 1.8550 0.6000 1.9450 1.4900 ;
      RECT 1.7500 0.5100 1.9450 0.6000 ;
      RECT 0.2400 0.9750 0.3300 1.0800 ;
      RECT 1.2300 1.1700 1.3200 1.4900 ;
      RECT 0.2400 1.0800 1.3200 1.1700 ;
  END
END NOR2B_X3M_A12TH

MACRO NOR2B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5600 ;
        RECT 0.5950 0.3200 0.6950 0.5600 ;
        RECT 1.1200 0.3200 1.2200 0.5950 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.6500 0.9600 0.7500 ;
        RECT 0.0450 0.7500 0.1450 1.4650 ;
        RECT 0.3350 0.5200 0.4350 0.6500 ;
        RECT 0.8600 0.5000 0.9600 0.6500 ;
        RECT 0.0450 1.4650 1.6050 1.5650 ;
        RECT 0.5900 1.5650 0.6800 1.8950 ;
        RECT 1.5050 1.5650 1.6050 1.9200 ;
    END
    ANTENNADIFFAREA 0.66775 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9250 1.0500 1.2550 1.1500 ;
        RECT 1.1650 1.1500 1.2550 1.2800 ;
        RECT 0.9250 1.1500 1.0150 1.2500 ;
        RECT 1.1650 1.2800 1.9250 1.3700 ;
        RECT 0.2350 1.2500 1.0150 1.3400 ;
        RECT 1.8350 0.9350 1.9250 1.2800 ;
        RECT 0.2350 0.9750 0.3250 1.2500 ;
        RECT 1.7950 0.7650 1.9250 0.9350 ;
    END
    ANTENNAGATEAREA 0.3084 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 1.0450 1.7700 1.1450 2.0800 ;
        RECT 1.9650 1.7700 2.0650 2.0800 ;
    END
  END VDD

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.8800 2.1500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END AN
  OBS
    LAYER M1 ;
      RECT 2.2300 1.5850 2.3300 1.9550 ;
      RECT 2.2400 0.7650 2.3300 1.5850 ;
      RECT 2.1850 0.6600 2.3300 0.7650 ;
      RECT 1.3650 0.5700 2.3300 0.6600 ;
      RECT 1.3650 1.0800 1.7450 1.1700 ;
      RECT 1.3650 0.6600 1.4550 0.8500 ;
      RECT 0.7450 0.8500 1.4550 0.9400 ;
      RECT 1.3650 0.9400 1.4550 1.0800 ;
      RECT 0.7450 0.9400 0.8350 1.0400 ;
      RECT 0.4550 1.0400 0.8350 1.1300 ;
  END
END NOR2B_X4M_A12TH

MACRO NOR2B_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.9450 0.3200 1.0450 0.6250 ;
        RECT 1.4650 0.3200 1.5650 0.6250 ;
        RECT 1.9850 0.3200 2.0850 0.6250 ;
        RECT 2.5050 0.3200 2.6050 0.6250 ;
        RECT 2.9050 0.3200 3.0050 0.6250 ;
        RECT 3.4250 0.3200 3.5250 0.6250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8350 1.0500 1.2250 1.1500 ;
        RECT 1.1250 1.0050 1.2250 1.0500 ;
        RECT 1.1250 0.9150 2.8450 1.0050 ;
        RECT 1.8550 1.0050 2.2250 1.1500 ;
        RECT 2.7550 0.7450 2.8450 0.9150 ;
    END
    ANTENNAGATEAREA 0.4626 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1350 1.0500 3.5550 1.1500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.4500 2.5450 1.5500 ;
        RECT 0.5350 1.5500 0.6350 1.8550 ;
        RECT 1.4650 1.5500 1.5650 1.8550 ;
        RECT 2.4450 1.5500 2.5450 1.8550 ;
        RECT 0.2450 0.8250 0.3450 1.4500 ;
        RECT 0.2450 0.7350 2.3450 0.8250 ;
        RECT 1.2050 0.4300 1.3050 0.7350 ;
        RECT 1.7250 0.4300 1.8250 0.7350 ;
        RECT 2.2450 0.4300 2.3450 0.7350 ;
    END
    ANTENNADIFFAREA 0.996 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.0750 1.7900 0.1750 2.0800 ;
        RECT 0.9950 1.7900 1.0950 2.0800 ;
        RECT 1.9850 1.7900 2.0850 2.0800 ;
        RECT 2.9050 1.4700 3.0050 2.0800 ;
        RECT 3.4250 1.4700 3.5250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4350 1.0000 0.5250 1.2400 ;
      RECT 0.4350 1.2400 3.2650 1.3300 ;
      RECT 2.9350 0.8700 3.2600 0.9600 ;
      RECT 2.9350 0.9600 3.0250 1.2400 ;
      RECT 3.1650 1.3300 3.2650 1.6600 ;
      RECT 3.1700 0.4350 3.2600 0.8700 ;
      RECT 1.3350 1.0950 1.7050 1.3300 ;
      RECT 2.3150 1.0950 2.6850 1.3300 ;
  END
END NOR2B_X6M_A12TH

MACRO NOR2B_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5800 ;
        RECT 0.5950 0.3200 0.6950 0.5800 ;
        RECT 1.1150 0.3200 1.2150 0.5800 ;
        RECT 1.6350 0.3200 1.7350 0.5800 ;
        RECT 2.1550 0.3200 2.2550 0.5800 ;
        RECT 4.1050 0.3200 4.2050 0.6100 ;
        RECT 4.6250 0.3200 4.7250 0.6100 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9800 1.0500 1.3500 1.1800 ;
        RECT 0.9800 1.1800 1.0700 1.2500 ;
        RECT 1.2600 1.1800 1.3500 1.2500 ;
        RECT 0.2350 1.2500 1.0700 1.3500 ;
        RECT 1.2600 1.2500 2.0550 1.3500 ;
        RECT 0.2350 1.0300 0.3250 1.2500 ;
        RECT 1.9650 1.1600 2.0550 1.2500 ;
        RECT 1.9650 1.0700 3.9350 1.1600 ;
        RECT 2.9750 1.1600 3.1850 1.2300 ;
        RECT 3.8450 1.1600 3.9350 1.2700 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2100 1.0500 4.6350 1.1550 ;
    END
    ANTENNAGATEAREA 0.1704 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.4500 3.5750 1.5500 ;
        RECT 0.5950 1.5500 0.6950 1.8600 ;
        RECT 1.6350 1.5500 1.7350 1.8600 ;
        RECT 2.5550 1.5500 2.6550 1.8600 ;
        RECT 3.4750 1.5500 3.5750 1.8600 ;
        RECT 0.0450 0.7800 0.1450 1.4500 ;
        RECT 0.0450 0.6800 1.9950 0.7800 ;
        RECT 0.3350 0.4100 0.4350 0.6800 ;
        RECT 0.8550 0.4100 0.9550 0.6800 ;
        RECT 1.3750 0.4100 1.4750 0.6800 ;
        RECT 1.8950 0.4100 1.9950 0.6800 ;
    END
    ANTENNADIFFAREA 1.328 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.0750 1.7900 0.1750 2.0800 ;
        RECT 1.1150 1.7900 1.2150 2.0800 ;
        RECT 2.0950 1.7900 2.1950 2.0800 ;
        RECT 3.0150 1.7900 3.1150 2.0800 ;
        RECT 4.0500 1.7050 4.1500 2.0800 ;
        RECT 4.6250 1.6750 4.7250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.3650 1.3550 4.4650 1.7000 ;
      RECT 4.0300 1.2650 4.4650 1.3550 ;
      RECT 4.0300 0.7600 4.4600 0.8500 ;
      RECT 4.3700 0.4550 4.4600 0.7600 ;
      RECT 4.0300 0.9600 4.1200 1.2650 ;
      RECT 1.7800 0.8700 4.1200 0.9600 ;
      RECT 4.0300 0.8500 4.1200 0.8700 ;
      RECT 0.7450 0.9600 0.8350 1.0600 ;
      RECT 0.4450 1.0600 0.8350 1.1500 ;
      RECT 1.4850 0.9600 1.5750 1.0700 ;
      RECT 0.7450 0.8700 1.5750 0.9600 ;
      RECT 1.7800 0.9600 1.8700 1.0700 ;
      RECT 1.4850 1.0700 1.8700 1.1600 ;
  END
END NOR2B_X8M_A12TH

MACRO NOR2XB_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4200 0.3200 0.5200 0.6000 ;
        RECT 0.9850 0.3200 1.1550 0.5050 ;
    END
  END VSS

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7500 0.3500 1.1700 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0050 0.9500 1.4600 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7000 1.1500 1.6600 ;
        RECT 0.9750 1.6600 1.1500 1.9800 ;
        RECT 0.7500 0.6100 1.1500 0.7000 ;
        RECT 0.7500 0.4100 0.8500 0.6100 ;
    END
    ANTENNADIFFAREA 0.120325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3750 1.6900 0.5450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.5000 0.6700 1.5900 ;
      RECT 0.5800 1.0300 0.6700 1.5000 ;
      RECT 0.0550 0.4500 0.2500 0.5400 ;
      RECT 0.0550 1.5900 0.1850 1.7400 ;
      RECT 0.0550 0.5400 0.1450 1.5000 ;
  END
END NOR2XB_X0P5M_A12TH

MACRO NOR2XB_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4200 0.3200 0.5200 0.6250 ;
        RECT 1.0150 0.3200 1.1250 0.5400 ;
    END
  END VSS

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7500 0.3500 1.1800 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8950 0.9500 1.3200 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7500 1.1500 1.7000 ;
        RECT 0.9750 1.7000 1.1500 1.9900 ;
        RECT 0.7500 0.6500 1.1500 0.7500 ;
        RECT 0.7500 0.4200 0.8500 0.6500 ;
    END
    ANTENNADIFFAREA 0.171175 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4400 1.7650 0.5500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.4600 0.7200 1.5500 ;
      RECT 0.6300 0.9700 0.7200 1.4600 ;
      RECT 0.0550 0.4750 0.2500 0.5650 ;
      RECT 0.0550 1.5500 0.1850 1.7400 ;
      RECT 0.0550 0.5650 0.1450 1.4600 ;
  END
END NOR2XB_X0P7M_A12TH

MACRO NOR2XB_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4350 0.3200 0.5350 0.8200 ;
        RECT 0.9250 0.3200 1.0950 0.7200 ;
    END
  END VSS

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.1550 0.3500 1.5950 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.5600 ;
        RECT 0.9800 1.5600 1.1500 1.6600 ;
        RECT 0.6950 0.8500 1.1500 0.9500 ;
        RECT 0.9800 1.6600 1.0800 1.9600 ;
        RECT 0.6950 0.4200 0.7950 0.8500 ;
    END
    ANTENNADIFFAREA 0.2752 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.1500 0.7500 1.4500 ;
        RECT 0.6500 1.0500 0.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4000 1.8950 0.5700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.7050 0.5400 1.7950 ;
      RECT 0.4500 0.9450 0.5400 1.7050 ;
      RECT 0.0500 0.6600 0.2500 0.7500 ;
      RECT 0.0500 0.7500 0.1400 1.7050 ;
  END
END NOR2XB_X1M_A12TH

MACRO NOR2XB_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3600 0.3200 0.4700 0.5200 ;
        RECT 0.8800 0.3200 0.9900 0.5300 ;
        RECT 1.4000 0.3200 1.5100 0.5300 ;
    END
  END VSS

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7650 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0333 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7500 1.5500 1.4500 ;
        RECT 0.8850 1.4500 1.5500 1.5500 ;
        RECT 0.6250 0.6500 1.5500 0.7500 ;
        RECT 0.8850 1.5500 0.9850 1.9050 ;
        RECT 0.6250 0.4250 0.7250 0.6500 ;
        RECT 1.1450 0.4250 1.2450 0.6500 ;
    END
    ANTENNADIFFAREA 0.235 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.4050 1.7000 1.5050 2.0800 ;
        RECT 0.4050 1.6800 0.5050 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.2500 1.1800 1.3500 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0500 1.3350 1.1400 ;
      RECT 1.2350 0.9300 1.3350 1.0500 ;
      RECT 0.0550 0.4100 0.2500 0.5000 ;
      RECT 0.0550 1.3900 0.1700 1.6800 ;
      RECT 0.0550 0.5000 0.1450 1.3000 ;
      RECT 0.0550 1.3000 0.5500 1.3900 ;
      RECT 0.4600 1.1400 0.5500 1.3000 ;
  END
END NOR2XB_X1P4M_A12TH

MACRO NOR2XB_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3300 0.3200 0.5000 0.6150 ;
        RECT 0.8800 0.3200 0.9900 0.4550 ;
        RECT 1.4000 0.3200 1.5100 0.4550 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7300 1.0500 1.1800 1.1500 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7650 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7500 1.5500 1.4500 ;
        RECT 0.8850 1.4500 1.5500 1.5500 ;
        RECT 0.6250 0.6500 1.5500 0.7500 ;
        RECT 0.8850 1.5500 0.9850 1.8900 ;
        RECT 0.6250 0.4350 0.7250 0.6500 ;
        RECT 1.1450 0.4300 1.2450 0.6500 ;
    END
    ANTENNADIFFAREA 0.332 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3550 1.7700 0.4550 2.0800 ;
        RECT 1.4050 1.7700 1.5050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5250 0.8600 1.3550 0.9500 ;
      RECT 0.0550 1.5000 0.6150 1.5900 ;
      RECT 0.5250 0.9500 0.6150 1.5000 ;
      RECT 0.0550 1.5900 0.1700 1.9700 ;
      RECT 0.0550 0.5550 0.1450 1.5000 ;
      RECT 0.0550 0.4650 0.2400 0.5550 ;
  END
END NOR2XB_X2M_A12TH

MACRO NOR2XB_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.5050 0.3200 0.6050 0.5600 ;
        RECT 1.0300 0.3200 1.1300 0.5600 ;
        RECT 1.5500 0.3200 1.6500 0.5950 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 1.3000 1.1500 ;
        RECT 0.2400 1.1500 0.3300 1.2500 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.7950 1.7500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0648 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7500 0.1500 1.4500 ;
        RECT 0.0500 1.4500 1.1300 1.5500 ;
        RECT 0.0500 0.6500 1.3900 0.7500 ;
        RECT 0.0500 1.5500 0.1700 1.9150 ;
        RECT 1.0300 1.5500 1.1300 1.9200 ;
        RECT 0.7700 0.5200 0.8700 0.6500 ;
        RECT 1.2900 0.5000 1.3900 0.6500 ;
    END
    ANTENNADIFFAREA 0.556425 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.5700 1.7700 0.6700 2.0800 ;
        RECT 1.5500 1.7700 1.6500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.8300 1.5700 1.9450 1.9550 ;
      RECT 1.4400 1.4800 1.9450 1.5700 ;
      RECT 1.8550 0.6000 1.9450 1.4800 ;
      RECT 1.7500 0.5100 1.9450 0.6000 ;
      RECT 1.4400 0.9600 1.5300 1.4800 ;
      RECT 0.4100 0.8500 1.5300 0.9600 ;
  END
END NOR2XB_X3M_A12TH

MACRO NOR2XB_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5600 ;
        RECT 0.5950 0.3200 0.6950 0.5600 ;
        RECT 1.1200 0.3200 1.2200 0.5950 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 1.0400 0.8350 1.1500 ;
        RECT 0.7450 0.9500 0.8350 1.0400 ;
        RECT 0.7450 0.8500 1.4550 0.9500 ;
        RECT 1.3650 0.9500 1.4550 1.0500 ;
        RECT 1.3650 1.0500 1.7450 1.1500 ;
    END
    ANTENNAGATEAREA 0.3084 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.8800 2.1500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.6500 0.9600 0.7500 ;
        RECT 0.0450 0.7500 0.1450 1.4650 ;
        RECT 0.3350 0.5200 0.4350 0.6500 ;
        RECT 0.8600 0.5000 0.9600 0.6500 ;
        RECT 0.0450 1.4650 1.6050 1.5650 ;
        RECT 0.5850 1.5650 0.6850 1.9200 ;
        RECT 1.5050 1.5650 1.6050 1.9200 ;
    END
    ANTENNADIFFAREA 0.66775 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 1.0450 1.7700 1.1450 2.0800 ;
        RECT 1.9650 1.7700 2.0650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2300 1.6650 2.3300 1.9550 ;
      RECT 1.8350 1.5750 2.3300 1.6650 ;
      RECT 2.2400 0.6750 2.3300 1.5750 ;
      RECT 2.1850 0.4800 2.3300 0.6750 ;
      RECT 1.8350 1.3550 1.9250 1.5750 ;
      RECT 0.2350 1.2650 1.9250 1.3550 ;
      RECT 1.8350 0.9150 1.9250 1.2650 ;
      RECT 1.7950 0.7450 1.9250 0.9150 ;
      RECT 1.0600 1.0500 1.1600 1.2650 ;
      RECT 0.2350 0.9750 0.3250 1.2650 ;
  END
END NOR2XB_X4M_A12TH

MACRO NOR2XB_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.9450 0.3200 1.0450 0.6250 ;
        RECT 1.4650 0.3200 1.5650 0.6250 ;
        RECT 1.9850 0.3200 2.0850 0.6250 ;
        RECT 2.5050 0.3200 2.6050 0.6250 ;
        RECT 2.9050 0.3200 3.0050 0.6250 ;
        RECT 3.4250 0.3200 3.5250 0.6250 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4350 1.2500 2.4150 1.3500 ;
        RECT 1.3350 1.2400 2.4150 1.2500 ;
        RECT 0.4350 1.0000 0.5250 1.2500 ;
        RECT 2.3150 1.1950 2.4150 1.2400 ;
        RECT 1.3350 1.0950 1.7050 1.2400 ;
        RECT 2.3150 1.0950 2.6850 1.1950 ;
    END
    ANTENNAGATEAREA 0.4626 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1350 1.0500 3.5550 1.1500 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.4500 2.5450 1.5500 ;
        RECT 0.5350 1.5500 0.6350 1.8550 ;
        RECT 1.4650 1.5500 1.5650 1.8550 ;
        RECT 2.4450 1.5500 2.5450 1.8550 ;
        RECT 0.2250 0.8250 0.3250 1.4500 ;
        RECT 0.2250 0.7350 2.3450 0.8250 ;
        RECT 1.2050 0.4300 1.3050 0.7350 ;
        RECT 1.7250 0.4300 1.8250 0.7350 ;
        RECT 2.2450 0.4300 2.3450 0.7350 ;
    END
    ANTENNADIFFAREA 0.996 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.0750 1.7900 0.1750 2.0800 ;
        RECT 0.9950 1.7900 1.0950 2.0800 ;
        RECT 1.9850 1.7900 2.0850 2.0800 ;
        RECT 2.9050 1.4700 3.0050 2.0800 ;
        RECT 3.4250 1.4700 3.5250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8350 1.0500 1.2250 1.1500 ;
      RECT 1.1250 1.0050 1.2250 1.0500 ;
      RECT 1.1250 0.9150 2.8950 1.0050 ;
      RECT 2.8050 1.2600 3.2650 1.3500 ;
      RECT 2.8050 0.7850 3.2600 0.8750 ;
      RECT 2.8050 0.8750 2.8950 0.9150 ;
      RECT 2.8050 1.0050 2.8950 1.2600 ;
      RECT 3.1650 1.3500 3.2650 1.6950 ;
      RECT 3.1700 0.4350 3.2600 0.7850 ;
      RECT 1.8550 0.9150 2.2250 1.1500 ;
  END
END NOR2XB_X6M_A12TH

MACRO NOR2XB_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5800 ;
        RECT 0.5950 0.3200 0.6950 0.5800 ;
        RECT 1.1150 0.3200 1.2150 0.5800 ;
        RECT 1.6350 0.3200 1.7350 0.5800 ;
        RECT 2.1550 0.3200 2.2550 0.5800 ;
        RECT 4.1050 0.3200 4.2050 0.6100 ;
        RECT 4.6250 0.3200 4.7250 0.6100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.0750 1.7900 0.1750 2.0800 ;
        RECT 1.1150 1.7900 1.2150 2.0800 ;
        RECT 2.0950 1.7900 2.1950 2.0800 ;
        RECT 3.0150 1.7900 3.1150 2.0800 ;
        RECT 4.0500 1.6750 4.1500 2.0800 ;
        RECT 4.6250 1.6750 4.7250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0500 0.8350 1.1500 ;
        RECT 0.7450 0.9600 0.8350 1.0500 ;
        RECT 0.7450 0.8700 1.5750 0.9600 ;
        RECT 1.4850 0.9600 1.5750 1.0700 ;
        RECT 1.4850 1.0700 1.8700 1.1600 ;
        RECT 1.7800 0.9600 1.8700 1.0700 ;
        RECT 1.7800 0.8700 3.5550 0.9600 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2100 1.0500 4.6350 1.1550 ;
    END
    ANTENNAGATEAREA 0.1704 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0550 1.4500 3.5750 1.5500 ;
        RECT 0.5950 1.5500 0.6950 1.8600 ;
        RECT 1.6350 1.5500 1.7350 1.8600 ;
        RECT 2.5550 1.5500 2.6550 1.8600 ;
        RECT 3.4750 1.5500 3.5750 1.8600 ;
        RECT 0.0550 0.7800 0.1450 1.4500 ;
        RECT 0.0550 0.6900 1.9950 0.7800 ;
        RECT 0.3350 0.4100 0.4350 0.6900 ;
        RECT 0.8550 0.4100 0.9550 0.6900 ;
        RECT 1.3750 0.4100 1.4750 0.6900 ;
        RECT 1.8950 0.4100 1.9950 0.6900 ;
    END
    ANTENNADIFFAREA 1.328 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 4.3650 1.3550 4.4650 1.6550 ;
      RECT 4.0300 1.2650 4.4650 1.3550 ;
      RECT 4.0300 0.7600 4.4600 0.8500 ;
      RECT 4.3700 0.4550 4.4600 0.7600 ;
      RECT 4.0300 1.1600 4.1200 1.2650 ;
      RECT 1.9650 1.0700 4.1200 1.1600 ;
      RECT 4.0300 0.8500 4.1200 1.0700 ;
      RECT 0.2350 1.0300 0.3250 1.2500 ;
      RECT 1.1100 1.0500 1.2100 1.2500 ;
      RECT 1.9650 1.1600 2.0550 1.2500 ;
      RECT 0.2350 1.2500 2.0550 1.3500 ;
      RECT 2.9750 1.1600 3.1850 1.2300 ;
  END
END NOR2XB_X8M_A12TH

MACRO NOR2_X0P5A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0850 0.3200 0.1950 0.7000 ;
        RECT 0.5750 0.3200 0.7450 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5250 0.1900 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8900 0.1600 1.3500 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0050 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8600 0.7500 1.5500 ;
        RECT 0.5500 1.5500 0.7500 1.6500 ;
        RECT 0.3500 0.7600 0.7500 0.8600 ;
        RECT 0.5500 1.6500 0.6500 1.9650 ;
        RECT 0.3500 0.5700 0.4500 0.7600 ;
    END
    ANTENNADIFFAREA 0.150275 ;
  END Y
END NOR2_X0P5A_A12TH

MACRO NOR2_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0650 0.3200 0.2350 0.6450 ;
        RECT 0.6150 0.3200 0.7250 0.7000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4350 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.8900 0.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8850 0.1500 1.5500 ;
        RECT 0.0500 1.5500 0.2150 1.9600 ;
        RECT 0.0500 0.7850 0.4600 0.8850 ;
        RECT 0.3600 0.4900 0.4600 0.7850 ;
    END
    ANTENNADIFFAREA 0.135 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6200 1.6700 0.7200 2.0800 ;
    END
  END VDD
END NOR2_X0P5B_A12TH

MACRO NOR2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0650 0.3200 0.2350 0.6450 ;
        RECT 0.6150 0.3200 0.7250 0.7000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.8900 0.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8850 0.1500 1.5500 ;
        RECT 0.0500 1.5500 0.2150 1.9600 ;
        RECT 0.0500 0.7850 0.4600 0.8850 ;
        RECT 0.3600 0.5100 0.4600 0.7850 ;
    END
    ANTENNADIFFAREA 0.116625 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6200 1.5250 0.7200 2.0800 ;
    END
  END VDD
END NOR2_X0P5M_A12TH

MACRO NOR2_X0P7A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.8650 ;
        RECT 0.6100 0.3200 0.7100 0.6750 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.1600 1.4100 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9000 0.7500 1.5500 ;
        RECT 0.5500 1.5500 0.7500 1.6500 ;
        RECT 0.3500 0.8000 0.7500 0.9000 ;
        RECT 0.5500 1.6500 0.6500 1.9600 ;
        RECT 0.3500 0.4750 0.4500 0.8000 ;
    END
    ANTENNADIFFAREA 0.213225 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5350 0.1900 2.0800 ;
    END
  END VDD
END NOR2_X0P7A_A12TH

MACRO NOR2_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7650 ;
        RECT 0.5750 0.3200 0.7450 0.6900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5350 0.1900 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.1600 1.4100 ;
    END
    ANTENNAGATEAREA 0.0477 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0477 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9000 0.7500 1.5500 ;
        RECT 0.5500 1.5500 0.7500 1.6500 ;
        RECT 0.3500 0.8000 0.7500 0.9000 ;
        RECT 0.5500 1.6500 0.6500 1.9600 ;
        RECT 0.3500 0.5550 0.4500 0.8000 ;
    END
    ANTENNADIFFAREA 0.162225 ;
  END Y
END NOR2_X0P7B_A12TH

MACRO NOR2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7950 ;
        RECT 0.5750 0.3200 0.7450 0.6900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5350 0.1900 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.1600 1.4100 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9000 0.7500 1.5500 ;
        RECT 0.5500 1.5500 0.7500 1.6500 ;
        RECT 0.3500 0.8000 0.7500 0.9000 ;
        RECT 0.5500 1.6500 0.6500 1.9600 ;
        RECT 0.3500 0.6400 0.4500 0.8000 ;
    END
    ANTENNADIFFAREA 0.185225 ;
  END Y
END NOR2_X0P7M_A12TH

MACRO NOR2_X1A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6900 ;
        RECT 0.6100 0.3200 0.7100 0.6900 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8950 0.3500 1.6500 ;
        RECT 0.2500 1.6500 0.7450 1.7500 ;
        RECT 0.2500 0.7950 0.4500 0.8950 ;
        RECT 0.5750 1.7500 0.7450 1.9700 ;
        RECT 0.3500 0.4200 0.4500 0.7950 ;
    END
    ANTENNADIFFAREA 0.27325 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0888 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5500 1.4550 ;
    END
    ANTENNAGATEAREA 0.0888 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0550 1.8700 0.2250 2.0800 ;
    END
  END VDD
END NOR2_X1A_A12TH

MACRO NAND4B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.7200 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0100 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7200 1.5500 1.7000 ;
        RECT 0.6450 1.7000 1.5500 1.8000 ;
        RECT 1.2100 0.6200 1.5500 0.7200 ;
        RECT 0.6450 1.8000 0.7450 1.9800 ;
        RECT 1.1700 1.8000 1.2600 1.9800 ;
        RECT 1.2100 0.4300 1.3800 0.6200 ;
    END
    ANTENNADIFFAREA 0.199375 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8950 1.2400 1.2800 1.3500 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.4500 1.1000 1.5700 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2400 0.5600 1.6350 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.9050 1.8900 1.0050 2.0800 ;
        RECT 1.4250 1.8900 1.5250 2.0800 ;
        RECT 0.3550 1.7950 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 0.8100 1.3600 0.9000 ;
      RECT 1.2700 0.9000 1.3600 1.0850 ;
      RECT 0.0500 1.8350 0.2250 1.9250 ;
      RECT 0.0500 0.9000 0.1400 1.8350 ;
      RECT 0.0500 0.6800 0.1400 0.8100 ;
      RECT 0.0500 0.5900 0.2250 0.6800 ;
  END
END NAND4B_X0P7M_A12TH

MACRO NAND4B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3300 0.3200 0.5000 0.9150 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.2800 0.7500 1.5050 ;
        RECT 0.6500 1.5050 0.9050 1.6500 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.4500 1.3300 1.6000 ;
        RECT 1.0500 1.2800 1.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.9050 2.0100 1.0050 2.0800 ;
        RECT 1.4250 2.0100 1.5250 2.0800 ;
        RECT 0.3550 1.8800 0.4550 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7200 1.5500 1.8200 ;
        RECT 0.6450 1.8200 1.5500 1.9200 ;
        RECT 1.2100 0.6200 1.5500 0.7200 ;
        RECT 0.6450 1.9200 0.7450 1.9900 ;
        RECT 1.1700 1.9200 1.2600 1.9900 ;
        RECT 1.2100 0.4300 1.3800 0.6200 ;
    END
    ANTENNADIFFAREA 0.28075 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2800 0.3500 1.7000 ;
    END
    ANTENNAGATEAREA 0.0219 ;
  END AN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2100 0.5600 1.6300 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.0550 1.0700 1.3400 1.1000 ;
      RECT 1.1200 1.1000 1.3400 1.1600 ;
      RECT 0.0550 1.0100 1.2100 1.0700 ;
      RECT 0.0550 1.9000 0.2250 1.9900 ;
      RECT 0.0550 1.1000 0.1450 1.9000 ;
      RECT 0.0550 0.8050 0.1850 1.0100 ;
  END
END NAND4B_X1M_A12TH

MACRO NAND4B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.5400 ;
        RECT 1.7550 0.3200 1.8550 0.7300 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3700 1.2500 1.4850 1.3550 ;
        RECT 0.3700 1.1600 0.4800 1.2500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0700 1.9500 1.4900 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6050 1.0500 1.3350 1.1600 ;
        RECT 1.1250 1.0250 1.3350 1.0500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.4500 1.6700 1.5700 ;
        RECT 1.4800 1.5700 1.6700 1.6450 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7500 0.1500 1.6700 ;
        RECT 0.0500 1.6700 1.0150 1.7700 ;
        RECT 0.0500 0.6500 1.0500 0.7500 ;
        RECT 0.3950 1.7700 0.4950 1.8900 ;
        RECT 0.9150 1.7700 1.0150 1.8900 ;
        RECT 0.8800 0.4100 1.0500 0.6500 ;
    END
    ANTENNADIFFAREA 0.317 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.1000 1.8800 0.2700 2.0800 ;
        RECT 0.6200 1.8800 0.7900 2.0800 ;
        RECT 1.1750 1.7700 1.2750 2.0800 ;
        RECT 1.7000 1.7500 1.8000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.9300 1.7050 2.1300 1.8050 ;
      RECT 2.0400 0.9300 2.1300 1.7050 ;
      RECT 0.7700 0.8400 2.1300 0.9300 ;
      RECT 2.0300 0.5850 2.1300 0.8400 ;
  END
END NAND4B_X1P4M_A12TH

MACRO NAND4B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6200 ;
        RECT 1.9550 0.3200 2.0550 0.8600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.6500 0.9900 1.7500 ;
        RECT 0.3000 1.7500 0.4700 1.9500 ;
        RECT 0.8200 1.7500 0.9900 1.9700 ;
        RECT 0.0450 0.8600 0.1450 1.6500 ;
        RECT 0.0450 0.7700 0.3550 0.8600 ;
        RECT 0.2650 0.7600 0.3550 0.7700 ;
        RECT 0.2650 0.6500 1.1800 0.7600 ;
        RECT 1.0100 0.4700 1.1800 0.6500 ;
    END
    ANTENNADIFFAREA 0.446 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.6500 1.8950 1.7500 ;
        RECT 1.2500 1.5500 1.3500 1.6500 ;
        RECT 0.2350 1.4500 1.3500 1.5500 ;
        RECT 0.2350 1.2350 0.3350 1.4500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.8500 1.7150 0.9500 ;
        RECT 0.4450 0.9500 0.5500 1.2000 ;
        RECT 1.6250 0.9500 1.7150 1.1900 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.5150 1.1500 ;
        RECT 0.7000 1.1500 0.8000 1.2900 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.1500 2.1500 1.6300 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END AN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.5600 1.8900 0.7300 2.0800 ;
        RECT 1.0800 1.8800 1.2500 2.0800 ;
        RECT 1.8450 1.8750 2.0200 2.0800 ;
        RECT 0.0750 1.8400 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1550 1.8900 2.3550 1.9900 ;
      RECT 2.2650 1.0400 2.3550 1.8900 ;
      RECT 1.8700 0.9500 2.3550 1.0400 ;
      RECT 2.2300 0.7900 2.3550 0.9500 ;
      RECT 1.8700 1.0400 1.9600 1.3350 ;
      RECT 1.0800 1.3350 1.9600 1.3400 ;
      RECT 1.4450 1.3400 1.9600 1.4250 ;
      RECT 1.0800 1.2400 1.5350 1.3350 ;
  END
END NAND4B_X2M_A12TH

MACRO NAND4B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.8550 ;
        RECT 1.3150 0.3200 1.4150 0.6300 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9600 0.3500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END AN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.2500 1.5700 1.3500 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.8250 1.1500 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9350 1.0500 3.0050 1.1500 ;
        RECT 1.9350 1.1500 2.0250 1.3000 ;
        RECT 2.5950 1.1500 3.0050 1.1950 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.6500 3.3550 1.7500 ;
        RECT 0.5600 1.7500 0.7300 1.9800 ;
        RECT 1.1200 1.7500 1.2100 1.9900 ;
        RECT 2.0000 1.7500 2.1700 1.9550 ;
        RECT 2.5200 1.7500 2.6900 1.9550 ;
        RECT 3.2650 0.9500 3.3550 1.6500 ;
        RECT 2.2350 0.8600 3.3550 0.9500 ;
        RECT 3.2300 0.5300 3.3550 0.8600 ;
    END
    ANTENNADIFFAREA 0.7172 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.8550 1.8450 0.9550 2.0800 ;
        RECT 1.3750 1.8450 1.4750 2.0800 ;
        RECT 1.7750 1.8450 1.8750 2.0800 ;
        RECT 2.3000 1.8450 2.3900 2.0800 ;
        RECT 2.8200 1.8450 2.9100 2.0800 ;
        RECT 0.3350 1.7500 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8600 0.7600 1.9200 0.8500 ;
      RECT 1.8300 0.5700 1.9200 0.7600 ;
      RECT 1.8300 0.4800 2.8900 0.5700 ;
      RECT 2.7200 0.5700 2.8900 0.7700 ;
      RECT 0.8600 0.4400 0.9500 0.7600 ;
      RECT 0.0500 1.4700 3.1550 1.5600 ;
      RECT 0.0500 1.5600 0.1700 1.8600 ;
      RECT 0.0500 0.8700 0.1400 1.4700 ;
      RECT 0.0500 0.6600 0.1700 0.8700 ;
  END
END NAND4B_X3M_A12TH

MACRO NAND4B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.8400 ;
        RECT 1.2550 0.3200 1.3550 0.6300 ;
        RECT 2.2300 0.3200 2.4000 0.5250 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9500 0.3500 1.3700 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END AN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 1.7250 1.8400 1.8250 2.0800 ;
        RECT 2.2450 1.8400 2.3450 2.0800 ;
        RECT 1.1750 1.7800 1.2750 2.0800 ;
        RECT 0.3350 1.7150 0.4350 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7600 1.0500 1.9900 1.1500 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1150 1.2500 2.2250 1.3500 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END D

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 1.2450 3.9500 1.7550 ;
        RECT 2.6950 1.7550 3.9500 1.8550 ;
        RECT 2.6950 1.2100 2.7950 1.7550 ;
    END
    ANTENNAGATEAREA 0.2724 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4150 1.6500 2.6050 1.7500 ;
        RECT 2.5050 1.1000 2.6050 1.6500 ;
        RECT 2.5050 1.0000 3.2450 1.1000 ;
        RECT 2.8850 1.1000 2.9850 1.4500 ;
        RECT 3.1450 0.9700 3.2450 1.0000 ;
        RECT 2.8850 1.4500 3.7300 1.5600 ;
        RECT 3.1450 0.8600 3.3550 0.9700 ;
        RECT 3.6300 1.1550 3.7300 1.4500 ;
        RECT 3.6300 1.0550 4.2250 1.1550 ;
        RECT 4.1250 1.1550 4.2250 1.4500 ;
        RECT 4.1250 1.4500 4.6350 1.5500 ;
        RECT 4.5350 0.7850 4.6350 1.4500 ;
        RECT 4.1800 0.6850 4.6350 0.7850 ;
    END
    ANTENNADIFFAREA 0.99275 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 3.4450 0.8750 4.4050 0.9650 ;
      RECT 4.3150 0.9650 4.4050 1.1900 ;
      RECT 0.0500 1.4600 2.4150 1.5500 ;
      RECT 2.3250 0.9100 2.4150 1.4600 ;
      RECT 0.0500 1.5500 0.1700 1.8900 ;
      RECT 0.0500 0.8600 0.1400 1.4600 ;
      RECT 0.0500 0.4900 0.1700 0.8600 ;
      RECT 2.3250 0.8200 2.9800 0.9100 ;
      RECT 2.8900 0.7500 2.9800 0.8200 ;
      RECT 2.8900 0.6600 3.5350 0.7500 ;
      RECT 3.4450 0.7500 3.5350 0.8750 ;
      RECT 3.4450 0.9650 3.5350 1.2400 ;
      RECT 3.1000 1.2400 3.5350 1.3500 ;
      RECT 2.7100 0.4800 4.8150 0.5700 ;
      RECT 4.7250 0.5700 4.8150 0.9100 ;
      RECT 1.7300 0.6400 2.8000 0.7300 ;
      RECT 2.7100 0.5700 2.8000 0.6400 ;
      RECT 3.7400 0.5700 3.9100 0.7850 ;
      RECT 0.8000 0.5200 0.8900 0.8600 ;
      RECT 0.8000 0.8600 1.8200 0.9500 ;
      RECT 1.7300 0.7300 1.8200 0.8600 ;
      RECT 1.7300 0.5200 1.8200 0.6400 ;
  END
END NAND4B_X4M_A12TH

MACRO NAND4XXXB_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.9000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8500 1.8900 1.0200 2.0800 ;
        RECT 1.3700 1.8900 1.5400 2.0800 ;
        RECT 0.3550 1.7900 0.4550 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.2400 1.0950 1.3500 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.4500 1.1000 1.5600 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END C

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0200 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END DN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0100 1.3500 1.1000 ;
        RECT 1.2500 1.1000 1.3500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.7000 ;
        RECT 0.6250 1.7000 1.5500 1.8000 ;
        RECT 1.1950 0.7600 1.5500 0.8600 ;
        RECT 0.6250 1.8000 0.7250 1.9800 ;
        RECT 1.1500 1.8000 1.2400 1.9800 ;
        RECT 1.1950 0.4800 1.2950 0.7600 ;
    END
    ANTENNADIFFAREA 0.139375 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0500 1.5000 0.5200 1.5900 ;
      RECT 0.4300 1.5900 0.5200 1.6700 ;
      RECT 0.0500 1.8500 0.2250 1.9400 ;
      RECT 0.0500 1.5900 0.1400 1.8500 ;
      RECT 0.0500 0.8700 0.1400 1.5000 ;
      RECT 0.0500 0.7800 0.2250 0.8700 ;
  END
END NAND4XXXB_X0P5M_A12TH

MACRO NAND4XXXB_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.8250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1850 1.1900 1.3500 ;
        RECT 0.8500 1.1000 0.9500 1.1850 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END B

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0100 0.3500 1.3700 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END DN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7000 1.5500 1.7000 ;
        RECT 0.6450 1.7000 1.5500 1.8000 ;
        RECT 1.2100 0.6000 1.5500 0.7000 ;
        RECT 0.6450 1.8000 0.7450 1.9900 ;
        RECT 1.1700 1.8000 1.2600 1.9900 ;
        RECT 1.2100 0.4100 1.3800 0.6000 ;
    END
    ANTENNADIFFAREA 0.199375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8700 1.8900 1.0400 2.0800 ;
        RECT 1.4250 1.8900 1.5250 2.0800 ;
        RECT 0.3550 1.7800 0.4550 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.4500 1.1000 1.5700 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1000 0.8100 1.3500 1.0450 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0500 1.5000 0.5550 1.5900 ;
      RECT 0.4650 1.5900 0.5550 1.6700 ;
      RECT 0.0500 1.8200 0.2250 1.9100 ;
      RECT 0.0500 1.5900 0.1400 1.8200 ;
      RECT 0.0500 0.7650 0.1400 1.5000 ;
      RECT 0.0500 0.6750 0.2250 0.7650 ;
  END
END NAND4XXXB_X0P7M_A12TH

MACRO NAND4XXXB_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3300 0.3200 0.5000 0.9150 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.3000 0.7550 1.5400 ;
        RECT 0.6500 1.5400 1.0250 1.6300 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0800 0.9500 1.3100 ;
        RECT 0.8500 1.3100 1.1050 1.4200 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7000 1.5500 1.7400 ;
        RECT 0.6450 1.7400 1.5500 1.8400 ;
        RECT 1.2100 0.6000 1.5500 0.7000 ;
        RECT 0.6450 1.8400 0.7450 1.9500 ;
        RECT 1.1700 1.8400 1.2600 1.9500 ;
        RECT 1.2100 0.4100 1.3800 0.6000 ;
    END
    ANTENNADIFFAREA 0.28075 ;
  END Y

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0500 0.3500 1.4700 ;
    END
    ANTENNAGATEAREA 0.0219 ;
  END DN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1500 1.0800 1.3500 1.1900 ;
        RECT 1.2450 0.8400 1.3500 1.0800 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8700 1.9600 1.0400 2.0800 ;
        RECT 1.4250 1.9450 1.5250 2.0800 ;
        RECT 0.3550 1.7650 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.5800 0.5600 1.6700 ;
      RECT 0.4600 1.5000 0.5600 1.5800 ;
      RECT 0.0500 1.8000 0.2250 1.8900 ;
      RECT 0.0500 1.6700 0.1400 1.8000 ;
      RECT 0.0500 0.9150 0.1400 1.5800 ;
      RECT 0.0500 0.8250 0.2250 0.9150 ;
  END
END NAND4XXXB_X1M_A12TH

MACRO NAND4XXXB_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6400 ;
        RECT 1.7550 0.3200 1.8550 0.7350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0550 1.9950 0.2250 2.0800 ;
        RECT 0.5750 1.8600 0.7450 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.7650 1.6700 1.8650 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.6500 1.0050 1.7500 ;
        RECT 0.3150 1.7500 0.4850 1.9650 ;
        RECT 0.8350 1.7500 1.0050 1.9650 ;
        RECT 0.0450 0.9500 0.1350 1.6500 ;
        RECT 0.0450 0.8500 0.3650 0.9500 ;
        RECT 0.2650 0.7500 0.3650 0.8500 ;
        RECT 0.2650 0.6500 1.0500 0.7500 ;
        RECT 0.8800 0.4200 1.0500 0.6500 ;
    END
    ANTENNADIFFAREA 0.317 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3100 1.0500 1.5550 1.1500 ;
        RECT 1.4550 1.1500 1.5550 1.2850 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 1.2500 1.3450 1.3500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7850 0.8500 1.2050 0.9500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END A

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8950 1.9650 1.3200 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END DN
  OBS
    LAYER M1 ;
      RECT 2.0300 1.5500 2.1450 1.7600 ;
      RECT 0.2250 1.4600 2.1450 1.5500 ;
      RECT 2.0550 0.7950 2.1450 1.4600 ;
      RECT 2.0300 0.5850 2.1450 0.7950 ;
      RECT 1.6450 0.8250 1.7350 1.4600 ;
      RECT 0.2250 1.3400 0.3150 1.4600 ;
  END
END NAND4XXXB_X1P4M_A12TH

MACRO NAND4XXXB_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6400 ;
        RECT 1.8900 0.3200 1.9900 0.6000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.6500 1.0100 1.7500 ;
        RECT 0.3100 1.7500 0.4800 1.9400 ;
        RECT 0.8400 1.7500 1.0100 1.9400 ;
        RECT 0.0450 0.9600 0.1450 1.6500 ;
        RECT 0.0450 0.8600 0.3650 0.9600 ;
        RECT 0.2650 0.7200 0.3650 0.8600 ;
        RECT 0.2650 0.6200 1.1600 0.7200 ;
        RECT 0.9900 0.4300 1.1600 0.6200 ;
    END
    ANTENNADIFFAREA 0.4533 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 0.8500 1.7150 0.9500 ;
        RECT 0.4550 0.9500 0.5550 1.2100 ;
        RECT 1.6250 0.9500 1.7150 1.3700 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9600 1.0400 1.3850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END A

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0100 2.1600 1.4300 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END DN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0750 1.9800 0.1750 2.0800 ;
        RECT 0.5700 1.8700 0.7400 2.0800 ;
        RECT 1.1300 1.7600 1.2350 2.0800 ;
        RECT 1.9150 1.7250 2.0850 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6550 1.2500 1.4700 1.3600 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END B
  OBS
    LAYER M1 ;
      RECT 2.2300 1.6350 2.3450 1.8700 ;
      RECT 1.7900 1.5500 2.3450 1.6350 ;
      RECT 0.2350 1.5450 2.3450 1.5500 ;
      RECT 2.2550 0.9250 2.3450 1.5450 ;
      RECT 2.2200 0.7150 2.3450 0.9250 ;
      RECT 0.2350 1.2200 0.3250 1.4600 ;
      RECT 0.2350 1.4600 1.8800 1.5450 ;
  END
END NAND4XXXB_X2M_A12TH

MACRO NAND4XXXB_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7550 ;
        RECT 1.2950 0.3200 1.3950 0.5600 ;
    END
  END VSS

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9300 0.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END DN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6550 1.0500 1.7500 1.1500 ;
        RECT 1.6500 1.1500 1.7500 1.2650 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8000 1.4500 2.9750 1.5500 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0650 1.2450 3.1500 1.3500 ;
        RECT 3.0500 1.1400 3.1500 1.2450 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5550 1.6500 3.3500 1.7500 ;
        RECT 0.5550 1.7500 0.7300 1.9500 ;
        RECT 1.1150 1.7500 1.2150 1.9900 ;
        RECT 1.9250 1.7500 2.1050 1.9550 ;
        RECT 2.4450 1.7500 2.6250 1.9550 ;
        RECT 3.2550 1.0300 3.3500 1.6500 ;
        RECT 2.2300 0.9400 3.3500 1.0300 ;
        RECT 2.2300 0.7600 2.3200 0.9400 ;
        RECT 3.2300 0.5400 3.3500 0.9400 ;
    END
    ANTENNADIFFAREA 0.7172 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.8550 1.8400 0.9550 2.0800 ;
        RECT 1.3750 1.8400 1.4750 2.0800 ;
        RECT 1.7050 1.8400 1.8050 2.0800 ;
        RECT 2.2250 1.8400 2.3250 2.0800 ;
        RECT 2.7450 1.8400 2.8450 2.0800 ;
        RECT 0.3350 1.7500 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.4400 1.5600 1.4650 ;
      RECT 1.1200 1.3750 1.5600 1.4400 ;
      RECT 0.0500 1.4650 1.2100 1.5300 ;
      RECT 0.0500 1.5300 0.1700 1.8500 ;
      RECT 0.0500 0.8400 0.1400 1.4400 ;
      RECT 0.0500 0.6300 0.1850 0.8400 ;
      RECT 1.7600 0.4800 2.8100 0.5700 ;
      RECT 2.7200 0.5700 2.8100 0.8500 ;
      RECT 0.8000 0.7800 1.8500 0.8700 ;
      RECT 1.7600 0.5700 1.8500 0.7800 ;
      RECT 0.8000 0.4400 0.8900 0.7800 ;
  END
END NAND4XXXB_X3M_A12TH

MACRO NAND4XXXB_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.5700 ;
        RECT 0.7600 0.3200 0.8600 0.5700 ;
        RECT 1.2800 0.3200 1.3800 0.5900 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5000 1.4400 2.9750 1.5500 ;
    END
    ANTENNAGATEAREA 0.2718 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6900 1.4400 2.2050 1.5500 ;
    END
    ANTENNAGATEAREA 0.2718 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1000 4.1500 1.7000 ;
        RECT 0.9850 1.7000 4.1500 1.8000 ;
        RECT 3.3600 1.0000 4.1500 1.1000 ;
        RECT 0.9850 1.8000 1.1550 1.9900 ;
        RECT 1.5050 1.8000 1.6750 1.9900 ;
        RECT 2.0250 1.8000 2.1950 1.9900 ;
        RECT 2.5450 1.8000 2.7150 1.9900 ;
        RECT 3.0650 1.8000 3.2350 1.9900 ;
        RECT 3.5850 1.8000 3.7550 1.9900 ;
        RECT 3.3600 0.6900 3.4600 1.0000 ;
        RECT 3.8800 0.6900 3.9800 1.0000 ;
    END
    ANTENNADIFFAREA 0.966375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2850 1.4400 3.7550 1.5500 ;
    END
    ANTENNAGATEAREA 0.2718 ;
  END A

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 0.7200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END DN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 1.2800 1.9100 1.3800 2.0800 ;
        RECT 1.8000 1.9100 1.9000 2.0800 ;
        RECT 2.3200 1.9100 2.4200 2.0800 ;
        RECT 2.8400 1.9100 2.9400 2.0800 ;
        RECT 3.3600 1.9100 3.4600 2.0800 ;
        RECT 3.8800 1.9100 3.9800 2.0800 ;
        RECT 0.3500 1.7000 0.4500 2.0800 ;
        RECT 0.7600 1.6900 0.8600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5100 1.4000 1.5300 ;
      RECT 0.8100 1.4400 1.4000 1.5100 ;
      RECT 0.0950 1.6000 0.1850 1.9300 ;
      RECT 0.0550 0.4450 0.2250 0.6600 ;
      RECT 0.0950 1.5300 0.9000 1.6000 ;
      RECT 0.8100 0.7500 0.9000 1.4400 ;
      RECT 0.0550 0.6600 0.9000 0.7500 ;
      RECT 1.0250 1.0100 1.6350 1.1000 ;
      RECT 1.5450 0.5700 1.6350 1.0100 ;
      RECT 1.5450 0.4800 2.1550 0.5700 ;
      RECT 2.0650 0.5700 2.1550 0.8900 ;
      RECT 1.0250 0.6700 1.1150 1.0100 ;
      RECT 1.8050 1.0100 2.4150 1.1000 ;
      RECT 1.8050 0.6900 1.8950 1.0100 ;
      RECT 2.3250 0.5700 2.4150 1.0100 ;
      RECT 2.3250 0.4800 2.9350 0.5700 ;
      RECT 2.8450 0.5700 2.9350 0.8900 ;
      RECT 3.1050 0.4800 3.7150 0.5700 ;
      RECT 3.6250 0.5700 3.7150 0.8900 ;
      RECT 2.5850 1.0100 3.1950 1.1000 ;
      RECT 2.5850 0.6900 2.6750 1.0100 ;
      RECT 3.1050 0.5700 3.1950 1.0100 ;
  END
END NAND4XXXB_X4M_A12TH

MACRO NAND4_X0P5A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1600 0.3200 0.2500 0.6800 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.7700 0.3600 1.1600 ;
    END
    ANTENNAGATEAREA 0.0411 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2950 1.2500 0.7150 1.3500 ;
    END
    ANTENNAGATEAREA 0.0411 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8900 1.1500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0411 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.0500 0.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.0411 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.4500 ;
        RECT 0.3650 1.4500 1.3500 1.5500 ;
        RECT 1.0900 0.6000 1.3500 0.7000 ;
        RECT 0.3650 1.5500 0.4650 1.7600 ;
        RECT 0.8900 1.5500 0.9800 1.7600 ;
    END
    ANTENNADIFFAREA 0.198925 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1100 1.6400 0.2000 2.0800 ;
        RECT 0.6300 1.6400 0.7200 2.0800 ;
        RECT 1.1550 1.6400 1.2450 2.0800 ;
    END
  END VDD
END NAND4_X0P5A_A12TH

MACRO NAND4_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1600 0.3200 0.2500 0.6800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6950 1.3500 1.4500 ;
        RECT 0.3650 1.4500 1.3500 1.5500 ;
        RECT 1.0900 0.5950 1.3500 0.6950 ;
        RECT 0.3650 1.5500 0.4650 1.8200 ;
        RECT 0.8900 1.5500 0.9800 1.8200 ;
    END
    ANTENNADIFFAREA 0.150925 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.0500 0.9200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8850 1.1500 1.3300 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2950 1.2500 0.7150 1.3500 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.7950 0.3650 1.1500 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1100 1.6400 0.2000 2.0800 ;
        RECT 0.6300 1.6400 0.7200 2.0800 ;
        RECT 1.1550 1.6400 1.2450 2.0800 ;
    END
  END VDD
END NAND4_X0P5M_A12TH

MACRO NAND4_X0P7A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 1.1450 0.3200 1.2350 0.8650 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9800 1.5500 ;
        RECT 0.3650 1.5500 0.4550 1.9850 ;
        RECT 0.8800 1.5500 0.9800 1.9850 ;
        RECT 0.2500 0.9000 0.3500 1.4500 ;
        RECT 0.1000 0.8000 0.3500 0.9000 ;
        RECT 0.1000 0.4700 0.2000 0.8000 ;
    END
    ANTENNADIFFAREA 0.265375 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8900 0.5500 1.3150 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9750 1.1600 1.3650 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0900 1.6400 0.1800 2.0800 ;
        RECT 0.6250 1.6400 0.7150 2.0800 ;
        RECT 1.1450 1.6400 1.2350 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0850 0.1600 1.5250 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8100 0.9500 1.1500 ;
        RECT 0.7400 1.1500 0.9500 1.2400 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END C
END NAND4_X0P7A_A12TH

MACRO NAND4_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 1.1450 0.3200 1.2350 0.8350 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8050 0.9500 1.1250 ;
        RECT 0.7500 1.1250 0.9500 1.2150 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0850 0.1600 1.5150 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9800 1.5500 ;
        RECT 0.3650 1.5500 0.4550 1.8100 ;
        RECT 0.8800 1.5500 0.9800 1.8100 ;
        RECT 0.2500 0.9700 0.3500 1.4500 ;
        RECT 0.1000 0.8700 0.3500 0.9700 ;
        RECT 0.1000 0.5600 0.2000 0.8700 ;
    END
    ANTENNADIFFAREA 0.199375 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0000 1.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END D

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8950 0.5500 1.3150 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1050 1.6500 0.1950 2.0800 ;
        RECT 0.6250 1.6500 0.7150 2.0800 ;
        RECT 1.1450 1.6500 1.2350 2.0800 ;
    END
  END VDD
END NAND4_X0P7M_A12TH

MACRO NAND4_X1A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 1.1450 0.3200 1.2350 0.6100 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8500 0.9500 1.1300 ;
        RECT 0.7700 1.1300 0.9500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0850 0.1600 1.5150 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9800 1.5500 ;
        RECT 0.3650 1.5500 0.4550 1.9200 ;
        RECT 0.8800 1.5500 0.9800 1.9200 ;
        RECT 0.2500 0.9700 0.3500 1.4500 ;
        RECT 0.1000 0.8700 0.3500 0.9700 ;
        RECT 0.1000 0.5600 0.2000 0.8700 ;
    END
    ANTENNADIFFAREA 0.37475 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7950 1.1500 1.2950 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END D

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8950 0.5500 1.3150 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0900 1.7000 0.1800 2.0800 ;
        RECT 0.6250 1.7000 0.7150 2.0800 ;
        RECT 1.1450 1.7000 1.2350 2.0800 ;
    END
  END VDD
END NAND4_X1A_A12TH

MACRO NAND4_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 1.1450 0.3200 1.2350 0.6100 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8000 0.9500 1.1550 ;
        RECT 0.7200 1.1550 0.9500 1.2550 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8900 0.5500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9050 1.1500 1.3550 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0950 0.1600 1.5050 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1050 1.6800 0.1950 2.0800 ;
        RECT 0.6250 1.6800 0.7150 2.0800 ;
        RECT 1.1450 1.5100 1.2350 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9800 1.5500 ;
        RECT 0.3650 1.5500 0.4550 1.9200 ;
        RECT 0.8800 1.5500 0.9800 1.9200 ;
        RECT 0.2500 0.9700 0.3500 1.4500 ;
        RECT 0.1000 0.8700 0.3500 0.9700 ;
        RECT 0.1000 0.5600 0.2000 0.8700 ;
    END
    ANTENNADIFFAREA 0.28075 ;
  END Y
END NAND4_X1M_A12TH

MACRO NAND4_X1P4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0650 0.3200 0.2350 0.5400 ;
        RECT 2.0000 0.3200 2.1000 0.6400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0750 1.9650 0.1750 2.0800 ;
        RECT 0.6200 1.8750 0.7900 2.0800 ;
        RECT 1.3250 1.7400 1.4250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9100 0.8400 1.4000 0.9500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.5550 1.1600 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.2500 1.7650 1.3500 ;
        RECT 1.6650 1.1050 1.7650 1.2500 ;
        RECT 0.4600 1.0050 0.5600 1.2500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.4500 1.9950 1.5500 ;
        RECT 1.8950 1.3050 1.9950 1.4500 ;
        RECT 0.2400 1.0050 0.3400 1.4500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6500 1.1550 0.7500 ;
        RECT 0.0500 0.7500 0.1500 1.6500 ;
        RECT 0.9850 0.4100 1.1550 0.6500 ;
        RECT 0.0500 1.6500 1.1050 1.7500 ;
        RECT 0.3050 1.7500 0.4750 1.9650 ;
        RECT 0.9350 1.7500 1.1050 1.9650 ;
    END
    ANTENNADIFFAREA 0.53825 ;
  END Y
END NAND4_X1P4A_A12TH

MACRO NAND4_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.4100 ;
        RECT 1.9950 0.3200 2.0950 0.6250 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.4500 1.9800 1.5500 ;
        RECT 0.2600 1.3500 0.3600 1.4500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 0.8500 1.7600 0.9500 ;
        RECT 0.4900 0.9500 0.5900 1.1800 ;
        RECT 1.6600 0.9500 1.7600 1.0900 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.2500 1.5250 1.3500 ;
        RECT 1.4350 1.1750 1.5250 1.2500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7250 1.0500 1.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6500 1.0950 1.7500 ;
        RECT 0.3000 1.7500 0.4700 1.9650 ;
        RECT 0.9250 1.7500 1.0950 1.9650 ;
        RECT 0.0500 0.7500 0.1500 1.6500 ;
        RECT 0.0500 0.6500 1.2100 0.7500 ;
        RECT 1.0400 0.4200 1.2100 0.6500 ;
    END
    ANTENNADIFFAREA 0.3586 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0750 1.9650 0.1750 2.0800 ;
        RECT 0.5800 1.8600 0.7500 2.0800 ;
        RECT 1.2600 1.7350 1.3600 2.0800 ;
    END
  END VDD
END NAND4_X1P4M_A12TH

MACRO NAND4_X2A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6300 ;
        RECT 2.2050 0.3200 2.2950 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9800 1.2500 1.4150 1.3500 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.0500 1.6250 1.1500 ;
        RECT 0.7700 1.1500 0.8700 1.2850 ;
        RECT 1.5250 1.1500 1.6250 1.2950 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.6500 ;
        RECT 0.3200 1.6500 2.3500 1.7500 ;
        RECT 1.9900 0.8500 2.3500 0.9500 ;
        RECT 0.3200 1.7500 0.4900 1.9800 ;
        RECT 0.8500 1.7500 1.0200 1.9750 ;
        RECT 1.3850 1.7500 1.5550 1.9750 ;
        RECT 1.9050 1.7500 2.0750 1.9750 ;
        RECT 1.9900 0.7500 2.0900 0.8500 ;
        RECT 1.1100 0.6500 2.0900 0.7500 ;
        RECT 1.1100 0.4300 1.2800 0.6500 ;
    END
    ANTENNADIFFAREA 0.6537 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2100 0.3500 1.4500 ;
        RECT 0.2500 1.4500 2.1500 1.5500 ;
        RECT 2.0500 1.2000 2.1500 1.4500 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5150 0.8500 1.8850 0.9500 ;
        RECT 0.5150 0.9500 0.6150 1.3050 ;
        RECT 1.7850 0.9500 1.8850 1.2600 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.6200 1.9100 0.7100 2.0800 ;
        RECT 1.1600 1.9100 1.2500 2.0800 ;
        RECT 1.6850 1.9100 1.7750 2.0800 ;
        RECT 2.2050 1.9100 2.2950 2.0800 ;
        RECT 0.0850 1.6850 0.1750 2.0800 ;
    END
  END VDD
END NAND4_X2A_A12TH

MACRO NAND4_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5600 ;
        RECT 1.9900 0.3200 2.0900 0.6400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0750 1.8400 0.1750 2.0800 ;
        RECT 0.6250 1.8400 0.7250 2.0800 ;
        RECT 1.1650 1.7700 1.2650 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.4500 1.9800 1.5500 ;
        RECT 0.2400 1.1400 0.3400 1.4500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4700 0.8500 1.7350 0.9500 ;
        RECT 0.4700 0.9500 0.5700 1.3450 ;
        RECT 1.6350 0.9500 1.7350 1.2750 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6850 1.2500 1.5150 1.3500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8750 1.0400 1.3000 1.1500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6500 1.0200 1.7500 ;
        RECT 0.3200 1.7500 0.4900 1.9600 ;
        RECT 0.8500 1.7500 1.0200 1.9650 ;
        RECT 0.0500 0.7500 0.1500 1.6500 ;
        RECT 0.0500 0.6500 1.1800 0.7500 ;
        RECT 1.0100 0.4350 1.1800 0.6500 ;
    END
    ANTENNADIFFAREA 0.4679 ;
  END Y
END NAND4_X2M_A12TH

MACRO NAND4_X3A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6300 ;
        RECT 0.6150 0.3200 0.7050 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8350 1.2500 2.3450 1.3500 ;
    END
    ANTENNAGATEAREA 0.2466 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.2500 0.8000 1.3500 ;
    END
    ANTENNAGATEAREA 0.2466 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0600 1.2500 1.5700 1.3500 ;
    END
    ANTENNAGATEAREA 0.2466 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6150 1.2500 3.1250 1.3500 ;
    END
    ANTENNAGATEAREA 0.2466 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0950 1.6450 0.1850 2.0800 ;
        RECT 0.6150 1.6450 0.7050 2.0800 ;
        RECT 1.1350 1.6450 1.2250 2.0800 ;
        RECT 1.6550 1.6450 1.7450 2.0800 ;
        RECT 2.1750 1.6450 2.2650 2.0800 ;
        RECT 2.6950 1.6450 2.7850 2.0800 ;
        RECT 3.2150 1.6450 3.3050 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.1500 3.3500 1.4500 ;
        RECT 0.3500 1.4500 3.3500 1.5500 ;
        RECT 2.6900 1.0500 3.3500 1.1500 ;
        RECT 0.3500 1.5500 0.4500 1.8900 ;
        RECT 0.8700 1.5500 0.9700 1.8900 ;
        RECT 1.3900 1.5500 1.4900 1.8900 ;
        RECT 1.9100 1.5500 2.0100 1.8900 ;
        RECT 2.4300 1.5500 2.5300 1.8900 ;
        RECT 2.9500 1.5500 3.0500 1.8900 ;
        RECT 2.6900 0.7600 2.7900 1.0500 ;
        RECT 3.2100 0.5400 3.3100 1.0500 ;
    END
    ANTENNADIFFAREA 0.9972 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.6550 0.8200 2.2650 0.9100 ;
      RECT 2.1750 0.6950 2.2650 0.8200 ;
      RECT 1.6550 0.5700 1.7450 0.8200 ;
      RECT 1.1350 0.4800 1.7450 0.5700 ;
      RECT 1.1350 0.5700 1.2250 0.6900 ;
      RECT 1.9150 0.4850 3.0450 0.5750 ;
      RECT 2.9550 0.5750 3.0450 0.9150 ;
      RECT 1.9150 0.5750 2.0050 0.7000 ;
      RECT 2.4350 0.5750 2.5250 0.9150 ;
      RECT 0.3550 0.8200 1.4850 0.9100 ;
      RECT 1.3950 0.6950 1.4850 0.8200 ;
      RECT 0.8750 0.4700 0.9650 0.8200 ;
      RECT 0.3550 0.4800 0.4450 0.8200 ;
  END
END NAND4_X3A_A12TH

MACRO NAND4_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 1.9600 0.3200 2.0600 0.6350 ;
        RECT 2.8950 0.3200 2.9950 0.6350 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4350 1.2500 1.3550 1.3500 ;
        RECT 1.2550 1.3500 1.3550 1.5000 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.8500 1.0900 0.9500 ;
        RECT 0.9900 0.9500 1.0900 1.0450 ;
        RECT 0.2450 0.9500 0.3450 1.2600 ;
        RECT 0.9900 1.0450 1.2550 1.1450 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7900 1.0500 2.9350 1.1500 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6500 2.8350 1.7500 ;
        RECT 0.5400 1.7500 0.7100 1.9850 ;
        RECT 1.0600 1.7500 1.2300 1.9850 ;
        RECT 2.1250 1.7500 2.2950 1.9850 ;
        RECT 2.6650 1.7500 2.8350 1.9850 ;
        RECT 1.4500 0.7600 1.5500 1.6500 ;
        RECT 0.0500 0.7400 0.1500 1.6500 ;
        RECT 0.9550 0.6600 1.5500 0.7600 ;
        RECT 0.0500 0.5300 0.2100 0.7400 ;
    END
    ANTENNADIFFAREA 0.75295 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6650 1.4500 2.6850 1.5500 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.2600 1.8550 0.4300 2.0800 ;
        RECT 0.8000 1.8550 0.9700 2.0800 ;
        RECT 1.3450 1.8550 1.5150 2.0800 ;
        RECT 1.8500 1.8550 2.0250 2.0800 ;
        RECT 2.3850 1.8550 2.5550 2.0800 ;
        RECT 2.9600 1.8550 3.1300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.7150 0.7400 2.5150 0.8300 ;
      RECT 2.4250 0.4200 2.5150 0.7400 ;
      RECT 1.7150 0.5700 1.8050 0.7400 ;
      RECT 0.5200 0.4800 1.8050 0.5700 ;
  END
END NAND4_X3M_A12TH

MACRO NAND4_X4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 2.2000 0.3200 2.3700 0.5200 ;
        RECT 3.1200 0.3200 3.2900 0.5200 ;
        RECT 4.1950 0.3200 4.2950 0.6300 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3400 1.2500 4.1900 1.3500 ;
        RECT 3.0150 1.1700 3.3950 1.2500 ;
        RECT 4.0900 1.0750 4.1900 1.2500 ;
        RECT 2.3400 1.0450 2.4400 1.2500 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8500 1.5200 0.9500 ;
        RECT 0.6500 0.9500 0.7500 1.0550 ;
        RECT 1.4200 0.9500 1.5200 1.0550 ;
        RECT 0.4450 1.0550 0.7500 1.1550 ;
        RECT 1.4200 1.0550 1.7000 1.1550 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.4500 4.0350 1.5500 ;
        RECT 0.7000 1.5500 0.8000 1.8800 ;
        RECT 1.2550 1.5500 1.3550 1.8800 ;
        RECT 1.7750 1.5500 1.8750 1.8800 ;
        RECT 2.8850 1.5500 2.9850 1.8800 ;
        RECT 3.4150 1.5500 3.5150 1.8800 ;
        RECT 3.9350 1.5500 4.0350 1.8850 ;
        RECT 2.0850 0.9450 2.1850 1.4500 ;
        RECT 1.7700 0.8450 2.1850 0.9450 ;
        RECT 1.7700 0.7600 1.8700 0.8450 ;
        RECT 0.4750 0.6600 1.8700 0.7600 ;
    END
    ANTENNADIFFAREA 1.332 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8050 0.8500 3.6900 0.9500 ;
        RECT 3.5900 0.9500 3.6900 1.0500 ;
        RECT 2.8050 0.9500 2.9050 1.0400 ;
        RECT 3.5900 1.0500 3.8850 1.1500 ;
        RECT 2.6450 1.0400 2.9050 1.1400 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1250 1.2500 1.9700 1.3500 ;
        RECT 0.8550 1.1700 1.2350 1.2500 ;
        RECT 1.8700 1.0850 1.9700 1.2500 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 0.4050 1.7700 0.5050 2.0800 ;
        RECT 0.9950 1.7700 1.0950 2.0800 ;
        RECT 1.5150 1.7700 1.6150 2.0800 ;
        RECT 2.0350 1.7700 2.1350 2.0800 ;
        RECT 2.5700 1.7700 2.6700 2.0800 ;
        RECT 3.1550 1.7700 3.2550 2.0800 ;
        RECT 3.6750 1.7700 3.7750 2.0800 ;
        RECT 4.1950 1.7700 4.2950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.9800 0.6550 3.8100 0.7450 ;
      RECT 3.6400 0.4350 3.8100 0.6550 ;
      RECT 0.0800 0.4800 2.0700 0.5700 ;
      RECT 1.9800 0.5700 2.0700 0.6550 ;
      RECT 0.0800 0.5700 0.1700 0.9100 ;
      RECT 2.6600 0.4300 2.8300 0.6550 ;
  END
END NAND4_X4A_A12TH

MACRO NAND3B_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.1000 0.3200 0.1900 0.6300 ;
        RECT 1.6600 0.3200 1.7500 0.6300 ;
        RECT 3.2200 0.3200 3.3100 0.6300 ;
        RECT 4.7800 0.3200 4.8700 0.6300 ;
        RECT 5.3750 0.3200 5.4650 0.9000 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5100 1.2500 4.4950 1.3500 ;
        RECT 0.5100 1.3500 0.6100 1.4700 ;
    END
    ANTENNAGATEAREA 0.4392 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.0500 4.7200 1.1500 ;
        RECT 0.2550 1.1500 0.3450 1.2800 ;
        RECT 4.6200 1.1500 4.7200 1.2600 ;
    END
    ANTENNAGATEAREA 0.4392 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0200 1.2500 5.4450 1.3500 ;
    END
    ANTENNAGATEAREA 0.123 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.6500 ;
        RECT 0.0500 1.6500 4.6500 1.7500 ;
        RECT 0.0500 0.8500 4.0900 0.9500 ;
        RECT 0.3200 1.7500 0.4900 1.9900 ;
        RECT 0.8400 1.7500 1.0100 1.9900 ;
        RECT 1.3600 1.7500 1.5300 1.9900 ;
        RECT 1.8800 1.7500 2.0500 1.9900 ;
        RECT 2.4000 1.7500 2.5700 1.9900 ;
        RECT 2.9200 1.7500 3.0900 1.9900 ;
        RECT 3.4400 1.7500 3.6100 1.9900 ;
        RECT 3.9600 1.7500 4.1300 1.9900 ;
        RECT 4.4800 1.7500 4.6500 1.9900 ;
        RECT 0.8800 0.5200 0.9700 0.8500 ;
        RECT 2.4400 0.5200 2.5300 0.8500 ;
        RECT 4.0000 0.5200 4.0900 0.8500 ;
    END
    ANTENNADIFFAREA 1.272 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.1000 1.9250 0.1900 2.0800 ;
        RECT 0.6150 1.9250 0.7150 2.0800 ;
        RECT 1.1350 1.9250 1.2350 2.0800 ;
        RECT 1.6550 1.9250 1.7550 2.0800 ;
        RECT 2.1750 1.9250 2.2750 2.0800 ;
        RECT 2.6950 1.9250 2.7950 2.0800 ;
        RECT 3.2150 1.9250 3.3150 2.0800 ;
        RECT 3.7350 1.9250 3.8350 2.0800 ;
        RECT 4.2550 1.9250 4.3550 2.0800 ;
        RECT 4.8400 1.7500 4.9300 2.0800 ;
        RECT 5.3750 1.7500 5.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 5.1150 1.5500 5.2050 1.9600 ;
      RECT 0.7250 1.4500 5.2050 1.5500 ;
      RECT 4.8100 1.0100 5.2050 1.1000 ;
      RECT 5.1150 0.5400 5.2050 1.0100 ;
      RECT 4.8100 1.1000 4.9000 1.4500 ;
  END
END NAND3B_X6M_A12TH

MACRO NAND3XXB_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3900 0.3200 0.5600 0.6500 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9100 1.8450 1.0800 2.0800 ;
        RECT 0.3600 1.7250 0.4600 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.0100 0.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0250 1.1500 1.4450 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 0.9800 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9000 1.3500 1.6450 ;
        RECT 0.6900 1.6450 1.3500 1.7550 ;
        RECT 1.2000 0.4850 1.3500 0.9000 ;
        RECT 0.6900 1.7550 0.7800 1.9500 ;
        RECT 1.2100 1.7550 1.3500 1.9450 ;
    END
    ANTENNADIFFAREA 0.15175 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5100 0.5800 1.6000 ;
      RECT 0.4900 0.8750 0.5800 1.5100 ;
      RECT 0.0450 0.7850 0.5800 0.8750 ;
      RECT 0.0950 1.6000 0.1850 1.9450 ;
  END
END NAND3XXB_X0P5M_A12TH

MACRO NAND3XXB_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3900 0.3200 0.5600 0.6650 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9100 1.8400 1.0800 2.0800 ;
        RECT 0.4250 1.7950 0.5250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0800 1.1500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END A

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 0.9850 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 0.9700 0.9500 1.3400 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8350 1.3500 1.6500 ;
        RECT 0.6900 1.6500 1.3500 1.7500 ;
        RECT 1.2000 0.4250 1.3500 0.8350 ;
        RECT 0.6900 1.7500 0.7800 1.8950 ;
        RECT 1.2100 1.7500 1.3500 1.8950 ;
    END
    ANTENNADIFFAREA 0.215375 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5100 0.5800 1.6000 ;
      RECT 0.4900 0.8750 0.5800 1.5100 ;
      RECT 0.0450 0.7850 0.5800 0.8750 ;
      RECT 0.0950 1.6000 0.1850 1.8950 ;
  END
END NAND3XXB_X0P7M_A12TH

MACRO NAND3XXB_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4250 0.3200 0.5250 0.6100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.4300 1.8600 0.5200 2.0800 ;
        RECT 0.9500 1.8600 1.0400 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.0150 0.9500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8500 1.3500 1.6500 ;
        RECT 0.6900 1.6500 1.3500 1.7500 ;
        RECT 1.2100 0.4400 1.3500 0.8500 ;
        RECT 0.6900 1.7500 0.7800 1.8950 ;
        RECT 1.2100 1.7500 1.3500 1.8950 ;
    END
    ANTENNADIFFAREA 0.3035 ;
  END Y

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.0550 0.3500 1.4650 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END CN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0800 1.1500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5850 0.5800 1.6750 ;
      RECT 0.4900 0.9200 0.5800 1.5850 ;
      RECT 0.0450 0.8300 0.5800 0.9200 ;
      RECT 0.0950 1.6750 0.1850 1.8300 ;
  END
END NAND3XXB_X1M_A12TH

MACRO NAND3XXB_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6500 ;
        RECT 1.3550 0.3200 1.4550 0.6500 ;
    END
  END VSS

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9000 1.7500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3700 1.0500 0.9500 1.1500 ;
        RECT 0.3700 1.1500 0.4700 1.2900 ;
        RECT 0.8400 1.1500 0.9500 1.3000 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 0.8500 0.9250 0.9500 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.4500 1.1500 1.5500 ;
        RECT 1.0500 0.7500 1.1500 1.4500 ;
        RECT 0.6800 0.6500 1.1500 0.7500 ;
        RECT 0.6800 0.4250 0.8500 0.6500 ;
    END
    ANTENNADIFFAREA 0.413 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.7050 2.0700 1.4900 2.0800 ;
        RECT 0.7050 1.9150 0.8750 2.0700 ;
        RECT 1.3200 1.9150 1.4900 2.0700 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1550 1.6550 1.9450 1.7450 ;
      RECT 1.8550 0.7000 1.9450 1.6550 ;
      RECT 1.6900 0.6100 1.9450 0.7000 ;
      RECT 1.2500 1.1050 1.3500 1.6550 ;
      RECT 0.1550 0.8250 0.2450 1.6550 ;
  END
END NAND3XXB_X1P4M_A12TH

MACRO NAND3XXB_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.4150 ;
        RECT 1.4350 0.3200 1.5350 0.5700 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5050 1.0500 0.9350 1.1800 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END A

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.0100 1.7600 1.4700 ;
    END
    ANTENNAGATEAREA 0.0423 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3050 1.4500 1.1650 1.5500 ;
        RECT 1.0500 1.0600 1.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 1.6500 1.3750 1.7500 ;
        RECT 0.6150 1.7500 0.7850 1.9400 ;
        RECT 1.1750 1.7500 1.2750 1.9800 ;
        RECT 1.2750 0.9500 1.3750 1.6500 ;
        RECT 0.6850 0.8500 1.3750 0.9500 ;
    END
    ANTENNADIFFAREA 0.5095 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.9150 1.8400 1.0150 2.0800 ;
        RECT 1.4350 1.8300 1.5350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.7700 1.6150 1.9450 1.8500 ;
      RECT 1.8550 0.8400 1.9450 1.6150 ;
      RECT 1.4650 0.7600 1.9450 0.8400 ;
      RECT 0.1850 0.6700 1.9450 0.7600 ;
      RECT 1.4650 0.8400 1.5550 1.2650 ;
      RECT 0.1850 0.7600 0.2750 1.2650 ;
  END
END NAND3XXB_X2M_A12TH

MACRO NAND3XXB_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.7300 0.3200 0.9000 0.5300 ;
        RECT 2.2100 0.3200 2.3100 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.4600 1.8500 0.6300 2.0800 ;
        RECT 1.0850 1.8500 1.2550 2.0800 ;
        RECT 1.6550 1.8500 1.8250 2.0800 ;
        RECT 2.2150 1.7550 2.3150 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0500 1.9500 1.1500 ;
        RECT 1.0500 1.1500 1.1500 1.2500 ;
        RECT 1.8500 1.1500 1.9500 1.3650 ;
        RECT 0.4100 1.2500 1.1500 1.3600 ;
        RECT 0.4100 1.0450 0.5100 1.2500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END B

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0450 2.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END CN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6500 2.0850 1.7500 ;
        RECT 0.7600 1.7500 0.9300 1.9550 ;
        RECT 1.3950 1.7500 1.5650 1.9550 ;
        RECT 1.9150 1.7500 2.0850 1.9550 ;
        RECT 0.0500 0.9700 0.1500 1.6500 ;
        RECT 0.0500 0.7500 0.2150 0.9700 ;
        RECT 0.0500 0.6500 1.5650 0.7500 ;
        RECT 0.0500 0.5400 0.2150 0.6500 ;
        RECT 1.3950 0.4500 1.5650 0.6500 ;
    END
    ANTENNADIFFAREA 0.70245 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.4500 1.3700 1.5500 ;
        RECT 1.2700 1.3500 1.3700 1.4500 ;
        RECT 1.2700 1.2500 1.6700 1.3500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END A
  OBS
    LAYER M1 ;
      RECT 2.5100 1.7100 2.6800 1.9700 ;
      RECT 2.5100 1.6200 2.7450 1.7100 ;
      RECT 2.6550 0.8550 2.7450 1.6200 ;
      RECT 0.8500 0.8450 2.7450 0.8550 ;
      RECT 2.1050 0.7650 2.7450 0.8450 ;
      RECT 2.5050 0.5150 2.6750 0.7650 ;
      RECT 0.8500 0.9350 0.9400 1.0300 ;
      RECT 0.6800 1.0300 0.9400 1.1300 ;
      RECT 0.8500 0.8550 2.2050 0.9350 ;
      RECT 2.1050 0.9350 2.2050 1.3050 ;
  END
END NAND3XXB_X3M_A12TH

MACRO NAND3XXB_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6300 ;
        RECT 1.3650 0.3200 1.5350 0.5300 ;
        RECT 2.9450 0.3200 3.1150 0.5300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 1.3600 1.8600 1.5300 2.0800 ;
        RECT 1.8850 1.8600 2.0550 2.0800 ;
        RECT 2.4200 1.8600 2.5900 2.0800 ;
        RECT 2.9800 1.8600 3.1500 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.2500 1.7000 1.3500 ;
        RECT 0.8400 1.0700 0.9400 1.2500 ;
        RECT 1.6000 0.9500 1.7000 1.2500 ;
        RECT 1.6000 0.8500 2.1500 0.9500 ;
        RECT 2.0500 0.9500 2.1500 1.0500 ;
        RECT 2.0500 1.0500 2.3450 1.1500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END A

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.0850 3.3500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0816 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7800 1.4500 2.6200 1.5500 ;
        RECT 1.8250 1.0450 1.9250 1.4500 ;
        RECT 2.5200 1.0450 2.6200 1.4500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5700 1.6500 2.8550 1.7500 ;
        RECT 1.6250 1.7500 1.7950 1.9650 ;
        RECT 2.1500 1.7500 2.3200 1.9650 ;
        RECT 2.6850 1.7500 2.8550 1.9650 ;
        RECT 2.7550 0.9350 2.8550 1.6500 ;
        RECT 0.5700 0.9150 0.6700 1.6500 ;
        RECT 2.4400 0.8350 2.8550 0.9350 ;
        RECT 0.5700 0.8150 0.9000 0.9150 ;
        RECT 2.4400 0.7600 2.5400 0.8350 ;
        RECT 2.1300 0.6600 2.5400 0.7600 ;
    END
    ANTENNADIFFAREA 0.848 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.1450 1.0900 0.4400 1.1800 ;
      RECT 0.3500 0.4800 1.1300 0.5700 ;
      RECT 0.3500 0.5700 0.4400 1.0900 ;
      RECT 1.0400 0.5700 1.1300 0.6700 ;
      RECT 1.0400 0.6700 1.7450 0.7600 ;
      RECT 1.3050 0.7600 1.4750 1.1450 ;
      RECT 1.6550 0.5700 1.7450 0.6700 ;
      RECT 1.6550 0.4800 2.7400 0.5700 ;
      RECT 2.6500 0.6300 3.0350 0.7200 ;
      RECT 2.6500 0.5700 2.7400 0.6300 ;
      RECT 2.9450 0.7200 3.0350 0.8050 ;
      RECT 2.9450 0.8950 3.0350 1.2150 ;
      RECT 2.9450 0.8050 3.5300 0.8950 ;
      RECT 3.3250 0.4650 3.4250 0.8050 ;
      RECT 3.4400 0.8950 3.5300 1.6650 ;
      RECT 3.2900 1.6650 3.5300 1.9650 ;
  END
END NAND3XXB_X4M_A12TH

MACRO NAND3XXB_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6450 ;
        RECT 1.6350 0.3200 1.7350 0.6250 ;
        RECT 3.1950 0.3200 3.2950 0.6500 ;
        RECT 4.8100 0.3200 4.9800 0.5050 ;
        RECT 5.4250 0.3200 5.5250 0.9400 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.2500 4.4050 1.3500 ;
        RECT 4.3150 1.1550 4.4050 1.2500 ;
    END
    ANTENNAGATEAREA 0.4392 ;
  END B

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0100 1.2500 5.4300 1.3500 ;
    END
    ANTENNAGATEAREA 0.123 ;
  END CN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.6850 4.6300 1.7500 ;
        RECT 0.3000 1.7500 0.4700 1.9900 ;
        RECT 0.8200 1.7500 0.9900 1.9900 ;
        RECT 1.3400 1.7500 1.5100 1.9900 ;
        RECT 1.8600 1.7500 2.0300 1.9900 ;
        RECT 2.3800 1.7500 2.5500 1.9900 ;
        RECT 2.9000 1.7500 3.0700 1.9900 ;
        RECT 3.4200 1.7500 3.5900 1.9900 ;
        RECT 3.9400 1.7500 4.1100 1.9900 ;
        RECT 4.4600 1.7500 4.6300 1.9900 ;
        RECT 0.0550 1.6500 4.6300 1.6850 ;
        RECT 0.0550 1.5950 0.4700 1.6500 ;
        RECT 4.5300 0.9550 4.6300 1.6500 ;
        RECT 0.0550 0.9500 0.1450 1.5950 ;
        RECT 3.9400 0.8500 4.6300 0.9550 ;
        RECT 0.0550 0.8500 2.5100 0.9500 ;
        RECT 3.9400 0.6650 4.1100 0.8500 ;
        RECT 0.0550 0.8400 0.9500 0.8500 ;
        RECT 2.4200 0.5200 2.5100 0.8500 ;
        RECT 0.8600 0.5200 0.9500 0.8400 ;
    END
    ANTENNADIFFAREA 1.272 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7250 1.4500 4.2050 1.5500 ;
    END
    ANTENNAGATEAREA 0.4392 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 3.6800 2.0100 3.8500 2.0800 ;
        RECT 4.2000 2.0100 4.3700 2.0800 ;
        RECT 0.5600 1.9950 0.7300 2.0800 ;
        RECT 1.0800 1.9950 1.2500 2.0800 ;
        RECT 1.6000 1.9950 1.7700 2.0800 ;
        RECT 2.1200 1.9950 2.2900 2.0800 ;
        RECT 2.6400 1.9950 2.8100 2.0800 ;
        RECT 3.1600 1.9950 3.3300 2.0800 ;
        RECT 4.8300 1.7800 4.9200 2.0800 ;
        RECT 5.4300 1.7800 5.5200 2.0800 ;
        RECT 0.0750 1.7750 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 5.1700 1.5800 5.2600 1.9700 ;
      RECT 4.7200 1.4900 5.2600 1.5800 ;
      RECT 4.7200 0.9950 5.2600 1.0850 ;
      RECT 5.1700 0.7150 5.2600 0.9950 ;
      RECT 4.5100 0.6250 5.2600 0.7150 ;
      RECT 4.7200 1.0850 4.8100 1.4900 ;
      RECT 0.2350 1.1600 0.3250 1.2800 ;
      RECT 4.5100 0.5750 4.6000 0.6250 ;
      RECT 3.5600 0.4850 4.6000 0.5750 ;
      RECT 3.5600 0.5750 3.6500 1.0700 ;
      RECT 0.2350 1.0700 3.6500 1.1600 ;
  END
END NAND3XXB_X6M_A12TH

MACRO NAND3_X0P5A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7200 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8850 0.7500 1.3050 ;
    END
    ANTENNAGATEAREA 0.0447 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.5500 1.1100 ;
        RECT 0.4050 1.1100 0.5500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0447 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8400 0.1600 1.2250 ;
    END
    ANTENNAGATEAREA 0.0447 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.7850 0.9500 1.4500 ;
        RECT 0.3050 1.4500 0.9500 1.5500 ;
        RECT 0.8150 0.4150 0.9500 0.7850 ;
        RECT 0.3050 1.5500 0.4050 1.8400 ;
        RECT 0.8200 1.5500 0.9500 1.6600 ;
    END
    ANTENNADIFFAREA 0.196975 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.0450 2.7200 ;
        RECT 0.0900 1.9700 0.1950 2.0800 ;
        RECT 0.5950 1.9700 0.6850 2.0800 ;
    END
  END VDD
END NAND3_X0P5A_A12TH

MACRO NAND3_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.8750 0.3200 0.9750 0.9150 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8950 0.1500 1.5000 ;
        RECT 0.0500 1.5000 0.7150 1.6000 ;
        RECT 0.0500 0.5100 0.1900 0.8950 ;
        RECT 0.0950 1.6000 0.1950 1.8400 ;
        RECT 0.6150 1.6000 0.7150 1.8400 ;
    END
    ANTENNADIFFAREA 0.1548 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3550 1.6900 0.4550 2.0800 ;
        RECT 0.8750 1.6900 0.9750 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.2100 0.9600 1.5900 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2900 0.7050 1.3900 ;
        RECT 0.4500 1.0950 0.5500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9700 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A
END NAND3_X0P5M_A12TH

MACRO NAND3_X0P7A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 1.0250 0.3200 1.1250 0.6550 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.8500 0.7500 1.2950 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9200 1.1500 1.1250 ;
        RECT 0.9250 1.1250 1.1500 1.2950 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7900 0.5500 1.4500 ;
        RECT 0.4500 1.4500 1.1250 1.5500 ;
        RECT 0.1900 0.6900 0.5500 0.7900 ;
        RECT 0.4500 1.5500 0.5600 1.9550 ;
        RECT 1.0250 1.5500 1.1250 1.9550 ;
        RECT 0.1900 0.4200 0.2800 0.6900 ;
    END
    ANTENNADIFFAREA 0.3035 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.1850 1.6400 0.2850 2.0800 ;
        RECT 0.7450 1.6400 0.8450 2.0800 ;
    END
  END VDD
END NAND3_X0P7A_A12TH

MACRO NAND3_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.9200 0.3200 1.0200 0.8100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9700 0.3500 1.3950 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9000 0.7500 1.2500 ;
        RECT 0.4950 1.2500 0.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9200 0.9500 1.3400 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8600 0.1500 1.5050 ;
        RECT 0.0500 1.5050 0.7600 1.6050 ;
        RECT 0.0500 0.7550 0.2250 0.8600 ;
        RECT 0.1400 1.6050 0.2400 1.9300 ;
        RECT 0.6600 1.6050 0.7600 1.9300 ;
        RECT 0.1250 0.4500 0.2250 0.7550 ;
    END
    ANTENNADIFFAREA 0.2495 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4000 1.6950 0.5000 2.0800 ;
        RECT 0.9200 1.5200 1.0200 2.0800 ;
    END
  END VDD
END NAND3_X0P7M_A12TH

MACRO NAND3_X1A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.9800 0.3200 1.0800 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9200 0.3550 1.3400 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.8250 1.1500 1.2800 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8100 0.1500 1.4500 ;
        RECT 0.0500 1.4500 0.8200 1.5500 ;
        RECT 0.0500 0.7100 0.3000 0.8100 ;
        RECT 0.2000 1.5500 0.3000 1.8250 ;
        RECT 0.7200 1.5500 0.8200 1.8800 ;
        RECT 0.2000 0.4400 0.3000 0.7100 ;
    END
    ANTENNADIFFAREA 0.44945 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9800 1.6800 1.0800 2.0800 ;
        RECT 0.4600 1.6700 0.5600 2.0800 ;
    END
  END VDD
END NAND3_X1A_A12TH

MACRO NAND3_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.8750 0.3200 0.9750 0.6000 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.0100 0.9600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9700 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3550 1.7550 0.4550 2.0800 ;
        RECT 0.8750 1.5350 0.9750 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2700 0.7050 1.3900 ;
        RECT 0.4500 1.0100 0.5500 1.2700 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8500 0.1500 1.5000 ;
        RECT 0.0500 1.5000 0.7150 1.6000 ;
        RECT 0.0500 0.7500 0.1950 0.8500 ;
        RECT 0.0950 1.6000 0.1950 1.9450 ;
        RECT 0.6150 1.6000 0.7150 1.9450 ;
        RECT 0.0950 0.4400 0.1950 0.7500 ;
    END
    ANTENNADIFFAREA 0.3096 ;
  END Y
END NAND3_X1M_A12TH

MACRO NAND3_X1P4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.6800 ;
        RECT 1.6550 0.3200 1.7550 0.6800 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.4500 1.6500 1.5500 ;
        RECT 1.5500 1.0750 1.6500 1.4500 ;
        RECT 0.2000 1.0200 0.3000 1.4500 ;
    END
    ANTENNAGATEAREA 0.1266 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 1.4000 1.3500 ;
        RECT 1.3000 1.0950 1.4000 1.2500 ;
        RECT 0.4500 0.9200 0.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.1266 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7350 1.0500 1.1750 1.1500 ;
    END
    ANTENNAGATEAREA 0.1266 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.6500 ;
        RECT 0.3200 1.6500 1.9500 1.7500 ;
        RECT 0.8750 0.8500 1.9500 0.9500 ;
        RECT 0.3200 1.7500 0.4900 1.9900 ;
        RECT 0.8400 1.7500 1.0100 1.9900 ;
        RECT 1.3600 1.7500 1.5300 1.9900 ;
        RECT 0.8750 0.4300 0.9750 0.8500 ;
    END
    ANTENNADIFFAREA 0.415 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.6150 1.8400 0.7150 2.0800 ;
        RECT 1.1350 1.8400 1.2350 2.0800 ;
        RECT 1.6550 1.8400 1.7550 2.0800 ;
        RECT 0.0950 1.7550 0.1950 2.0800 ;
    END
  END VDD
END NAND3_X1P4A_A12TH

MACRO NAND3_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6000 ;
        RECT 1.4300 0.3200 1.5200 0.6500 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.4500 1.4200 1.5500 ;
        RECT 1.3200 1.3300 1.4200 1.4500 ;
        RECT 0.2600 1.2500 0.3600 1.4500 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.2500 1.1750 1.3500 ;
        RECT 0.4850 1.1300 0.5950 1.2500 ;
        RECT 1.0850 1.1300 1.1750 1.2500 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.8500 1.0150 0.9950 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.6500 0.9200 0.7500 ;
        RECT 0.2500 0.7500 0.3500 1.0000 ;
        RECT 0.7500 0.4600 0.9200 0.6500 ;
        RECT 0.0500 1.0000 0.3500 1.1000 ;
        RECT 0.0500 1.1000 0.1500 1.6400 ;
        RECT 0.0500 1.6400 0.9900 1.7300 ;
        RECT 0.3350 1.7300 0.4350 1.9900 ;
        RECT 0.8200 1.7300 0.9900 1.9300 ;
    END
    ANTENNADIFFAREA 0.3522 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.0800 1.8200 0.1700 2.0800 ;
        RECT 0.6000 1.8200 0.6900 2.0800 ;
    END
  END VDD
END NAND3_X1P4M_A12TH

MACRO NAND3_X2A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.6300 ;
        RECT 1.6550 0.3200 1.7550 0.6300 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 1.6500 1.5500 ;
        RECT 0.2500 1.1000 0.3500 1.4500 ;
        RECT 1.5500 1.1000 1.6500 1.4500 ;
    END
    ANTENNAGATEAREA 0.1788 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5000 1.2500 1.3900 1.3500 ;
        RECT 0.5000 1.1000 0.6150 1.2500 ;
        RECT 1.2900 1.1000 1.3900 1.2500 ;
    END
    ANTENNAGATEAREA 0.1788 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7450 1.0500 1.1800 1.1500 ;
    END
    ANTENNAGATEAREA 0.1788 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.6500 ;
        RECT 0.3200 1.6500 1.9500 1.7500 ;
        RECT 0.8750 0.8500 1.9500 0.9500 ;
        RECT 0.3200 1.7500 0.4900 1.9900 ;
        RECT 0.8750 1.7500 0.9750 1.9900 ;
        RECT 1.3950 1.7500 1.4950 1.9900 ;
        RECT 0.8750 0.5200 0.9750 0.8500 ;
    END
    ANTENNADIFFAREA 0.586 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.5800 1.8500 0.7500 2.0800 ;
        RECT 1.1000 1.8500 1.2700 2.0800 ;
        RECT 1.6200 1.8500 1.7900 2.0800 ;
        RECT 0.0950 1.7400 0.1950 2.0800 ;
    END
  END VDD
END NAND3_X2A_A12TH

MACRO NAND3_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1800 0.5600 ;
        RECT 1.6050 0.3200 1.6950 0.6250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.0900 1.8400 0.1800 2.0800 ;
        RECT 0.6100 1.8400 0.7000 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.4500 1.6500 1.5500 ;
        RECT 0.2450 1.0300 0.3450 1.4500 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.2500 1.4150 1.3600 ;
        RECT 0.4950 1.0300 0.5950 1.2500 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7150 1.0500 1.1000 1.1600 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6500 1.0000 0.7500 ;
        RECT 0.0500 0.7500 0.1500 1.6500 ;
        RECT 0.8300 0.4400 1.0000 0.6500 ;
        RECT 0.0500 1.6500 1.0000 1.7400 ;
        RECT 0.3450 1.7400 0.4450 1.9900 ;
        RECT 0.8300 1.7400 1.0000 1.9400 ;
    END
    ANTENNADIFFAREA 0.478 ;
  END Y
END NAND3_X2M_A12TH

MACRO NAND3_X3A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6300 ;
        RECT 0.5950 0.3200 0.6950 0.6300 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0500 0.7200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2682 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9000 1.7500 1.3000 ;
        RECT 0.3350 1.3000 2.5150 1.4000 ;
        RECT 1.6500 0.8000 2.5100 0.9000 ;
        RECT 0.3350 1.4000 0.4350 1.7300 ;
        RECT 0.8550 1.4000 0.9550 1.7300 ;
        RECT 1.3750 1.4000 1.4750 1.7300 ;
        RECT 1.8950 1.4000 1.9950 1.7300 ;
        RECT 2.4150 1.4000 2.5150 1.7300 ;
        RECT 2.4200 0.4900 2.5100 0.8000 ;
    END
    ANTENNADIFFAREA 0.9684 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0800 1.0500 1.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2682 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8800 1.0500 2.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2682 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.0750 1.5800 0.1750 2.0800 ;
        RECT 0.5950 1.5800 0.6950 2.0800 ;
        RECT 1.1150 1.5800 1.2150 2.0800 ;
        RECT 1.6350 1.5800 1.7350 2.0800 ;
        RECT 2.1550 1.5800 2.2550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3350 0.8100 1.4750 0.9000 ;
      RECT 1.3750 0.6900 1.4750 0.8100 ;
      RECT 0.8550 0.4700 0.9550 0.8100 ;
      RECT 0.3350 0.4700 0.4350 0.8100 ;
      RECT 1.0600 0.4800 2.3100 0.5700 ;
  END
END NAND3_X3A_A12TH

MACRO NAND3_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6300 ;
        RECT 0.5950 0.3200 0.6950 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0800 1.0500 1.5250 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.0500 0.7200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9000 1.7500 1.2800 ;
        RECT 0.3350 1.2800 2.5150 1.3800 ;
        RECT 1.6500 0.8000 2.5150 0.9000 ;
        RECT 0.3350 1.3800 0.4350 1.8050 ;
        RECT 0.8550 1.3800 0.9550 1.8050 ;
        RECT 1.3750 1.3800 1.4750 1.8050 ;
        RECT 1.8950 1.3800 1.9950 1.8050 ;
        RECT 2.4150 1.3800 2.5150 1.8050 ;
        RECT 2.4150 0.4850 2.5150 0.8000 ;
    END
    ANTENNADIFFAREA 0.7092 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8700 1.0500 2.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.5950 1.4800 0.6950 2.0800 ;
        RECT 1.1150 1.4800 1.2150 2.0800 ;
        RECT 1.6350 1.4800 1.7350 2.0800 ;
        RECT 2.1550 1.4800 2.2550 2.0800 ;
        RECT 0.0750 1.3850 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3350 0.8100 1.4750 0.9000 ;
      RECT 1.3750 0.6900 1.4750 0.8100 ;
      RECT 0.8550 0.4800 0.9550 0.8100 ;
      RECT 0.3350 0.4900 0.4350 0.8100 ;
      RECT 1.0600 0.4800 2.3100 0.5700 ;
  END
END NAND3_X3M_A12TH

MACRO NAND3_X4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.6300 ;
        RECT 1.6200 0.3200 1.7900 0.5450 ;
        RECT 3.2150 0.3200 3.3150 0.6300 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 1.4500 3.1550 1.5500 ;
        RECT 1.7950 1.3500 1.8950 1.4500 ;
        RECT 3.0550 1.1050 3.1550 1.4500 ;
        RECT 1.5100 1.2500 1.8950 1.3500 ;
        RECT 1.5100 1.3500 1.6100 1.4500 ;
        RECT 0.2500 1.4500 1.6100 1.5500 ;
        RECT 0.2500 1.1100 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.3576 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.9500 3.3500 1.6400 ;
        RECT 0.3200 1.6400 3.3500 1.7400 ;
        RECT 2.4400 0.8500 3.3500 0.9500 ;
        RECT 0.3200 1.7400 0.4900 1.9900 ;
        RECT 0.8750 1.7400 0.9750 1.9900 ;
        RECT 1.3950 1.7400 1.4950 1.9900 ;
        RECT 1.9150 1.7400 2.0150 1.9900 ;
        RECT 2.4350 1.7400 2.5350 1.9900 ;
        RECT 2.9550 1.7400 3.0550 1.9900 ;
        RECT 2.4400 0.7500 2.5400 0.8500 ;
        RECT 0.8400 0.6500 2.5400 0.7500 ;
        RECT 2.4400 0.5200 2.5400 0.6500 ;
        RECT 0.8400 0.4400 1.0100 0.6500 ;
    END
    ANTENNADIFFAREA 1.172 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5100 1.2500 1.3950 1.3500 ;
        RECT 1.2950 1.1500 1.3950 1.2500 ;
        RECT 0.5100 1.1100 0.6100 1.2500 ;
        RECT 1.2950 1.0500 2.1200 1.1500 ;
        RECT 2.0200 1.1500 2.1200 1.2500 ;
        RECT 2.0200 1.2500 2.9000 1.3500 ;
        RECT 2.8000 1.1050 2.9000 1.2500 ;
    END
    ANTENNAGATEAREA 0.3576 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0550 0.8500 2.3500 0.9500 ;
        RECT 1.0550 0.9500 1.1550 1.0500 ;
        RECT 2.2500 0.9500 2.3500 1.0500 ;
        RECT 0.7250 1.0500 1.1550 1.1500 ;
        RECT 2.2500 1.0500 2.6650 1.1500 ;
    END
    ANTENNAGATEAREA 0.3576 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 3.1800 1.8600 3.3500 2.0800 ;
        RECT 0.6150 1.8300 0.7150 2.0800 ;
        RECT 1.1350 1.8300 1.2350 2.0800 ;
        RECT 1.6550 1.8300 1.7550 2.0800 ;
        RECT 2.1750 1.8300 2.2750 2.0800 ;
        RECT 2.6950 1.8300 2.7950 2.0800 ;
        RECT 0.0950 1.7500 0.1950 2.0800 ;
    END
  END VDD
END NAND3_X4A_A12TH

MACRO NAND3_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6300 ;
        RECT 1.6450 0.3200 1.7350 0.6300 ;
        RECT 3.2300 0.3200 3.3200 0.6300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.6500 ;
        RECT 0.0500 1.6500 3.3400 1.7500 ;
        RECT 0.0500 0.8500 0.9500 0.9500 ;
        RECT 0.3450 1.7500 0.4350 1.8950 ;
        RECT 0.8650 1.7500 0.9550 1.8950 ;
        RECT 1.3850 1.7500 1.4750 1.8950 ;
        RECT 1.9050 1.7500 1.9950 1.8950 ;
        RECT 2.4450 1.7500 2.5350 1.8950 ;
        RECT 2.9650 1.7500 3.0550 1.8950 ;
        RECT 3.2500 0.9500 3.3400 1.6500 ;
        RECT 0.8600 0.5200 0.9500 0.8500 ;
        RECT 2.4500 0.8500 3.3400 0.9500 ;
        RECT 2.4500 0.5200 2.5400 0.8500 ;
    END
    ANTENNADIFFAREA 0.8711 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 2.9050 1.3500 ;
        RECT 2.8150 1.1300 2.9050 1.2500 ;
        RECT 0.4500 1.0600 0.5400 1.2500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7200 1.0500 2.5850 1.1600 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 3.1400 1.5500 ;
        RECT 0.2500 1.3400 0.3600 1.4500 ;
        RECT 3.0350 1.2350 3.1400 1.4500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0750 1.9250 0.1850 2.0800 ;
        RECT 0.6050 1.9250 0.6950 2.0800 ;
        RECT 1.1250 1.9250 1.2150 2.0800 ;
        RECT 1.6450 1.9250 1.7350 2.0800 ;
        RECT 2.1650 1.9250 2.2550 2.0800 ;
        RECT 2.7050 1.9250 2.7950 2.0800 ;
        RECT 3.2250 1.9250 3.3150 2.0800 ;
    END
  END VDD
END NAND3_X4M_A12TH

MACRO NAND3_X6A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6400 ;
        RECT 0.8550 0.3200 0.9550 0.6400 ;
        RECT 1.3750 0.3200 1.4750 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 3.7450 1.7700 3.8450 2.0800 ;
        RECT 4.2650 1.7700 4.3650 2.0800 ;
        RECT 0.0750 1.7300 0.1750 2.0800 ;
        RECT 0.5950 1.7300 0.6950 2.0800 ;
        RECT 1.1150 1.7300 1.2150 2.0800 ;
        RECT 1.6500 1.6500 1.7500 2.0800 ;
        RECT 2.1700 1.6500 2.2700 2.0800 ;
        RECT 2.6900 1.6500 2.7900 2.0800 ;
        RECT 3.2250 1.6500 3.3250 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9000 1.2500 2.8550 1.3500 ;
    END
    ANTENNAGATEAREA 0.5364 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2000 1.0500 4.4300 1.1500 ;
    END
    ANTENNAGATEAREA 0.5364 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3350 1.4500 4.6250 1.5450 ;
        RECT 1.3750 1.5450 4.6250 1.5500 ;
        RECT 0.3350 1.5450 0.4350 1.8750 ;
        RECT 0.8550 1.5450 0.9550 1.8750 ;
        RECT 0.3350 1.4450 1.4750 1.4500 ;
        RECT 2.9650 0.9000 3.0650 1.4500 ;
        RECT 1.3750 1.5500 1.4750 1.8900 ;
        RECT 1.9100 1.5500 2.0100 1.8800 ;
        RECT 2.4300 1.5500 2.5300 1.8800 ;
        RECT 2.9450 1.5500 3.0650 1.8950 ;
        RECT 3.4850 1.5500 3.5850 1.8800 ;
        RECT 4.0050 1.5500 4.1050 1.8800 ;
        RECT 4.5250 1.5500 4.6250 1.8800 ;
        RECT 2.9650 0.8000 4.4200 0.9000 ;
    END
    ANTENNADIFFAREA 1.82675 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.0500 1.5150 1.1500 ;
    END
    ANTENNAGATEAREA 0.5364 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.0750 0.8100 2.8400 0.9000 ;
      RECT 1.6500 0.4700 1.7500 0.8100 ;
      RECT 0.0750 0.4700 0.1750 0.8100 ;
      RECT 0.5950 0.4700 0.6950 0.8100 ;
      RECT 1.1150 0.4700 1.2150 0.8100 ;
      RECT 4.5250 0.5700 4.6250 0.9100 ;
      RECT 1.8550 0.4800 4.6250 0.5700 ;
  END
END NAND3_X6A_A12TH

MACRO NAND3_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6400 ;
        RECT 0.8550 0.3200 0.9550 0.6400 ;
        RECT 1.3750 0.3200 1.4750 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 1.6500 1.6950 1.7500 2.0800 ;
        RECT 2.1350 1.6700 2.3050 2.0800 ;
        RECT 2.6550 1.6700 2.8250 2.0800 ;
        RECT 0.0750 1.4900 0.1750 2.0800 ;
        RECT 0.5950 1.4900 0.6950 2.0800 ;
        RECT 1.1150 1.4900 1.2150 2.0800 ;
        RECT 3.2250 1.4900 3.3250 2.0800 ;
        RECT 3.7450 1.4900 3.8450 2.0800 ;
        RECT 4.2650 1.4900 4.3650 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9000 1.2500 2.8550 1.3500 ;
    END
    ANTENNAGATEAREA 0.438 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2000 1.0500 4.4300 1.1500 ;
    END
    ANTENNAGATEAREA 0.4392 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3750 1.4500 3.0650 1.5500 ;
        RECT 1.3750 1.5500 1.4750 1.8700 ;
        RECT 1.9100 1.5500 2.0100 1.8800 ;
        RECT 2.4300 1.5500 2.5300 1.8800 ;
        RECT 2.9450 1.5500 3.0650 1.8800 ;
        RECT 1.3750 1.4000 1.4750 1.4500 ;
        RECT 2.9650 1.4000 3.0650 1.4500 ;
        RECT 0.3350 1.3000 1.4750 1.4000 ;
        RECT 2.9650 1.3000 4.6250 1.4000 ;
        RECT 0.3350 1.4000 0.4350 1.8700 ;
        RECT 0.8550 1.4000 0.9550 1.8700 ;
        RECT 3.4850 1.4000 3.5850 1.8700 ;
        RECT 4.0050 1.4000 4.1050 1.8700 ;
        RECT 4.5250 1.4000 4.6250 1.8700 ;
        RECT 2.9650 0.9000 3.0650 1.3000 ;
        RECT 2.9650 0.8000 4.4200 0.9000 ;
    END
    ANTENNADIFFAREA 1.31385 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.0500 1.5150 1.1500 ;
    END
    ANTENNAGATEAREA 0.4392 ;
  END C
  OBS
    LAYER M1 ;
      RECT 0.0750 0.8100 2.8400 0.9000 ;
      RECT 1.6500 0.4700 1.7500 0.8100 ;
      RECT 0.0750 0.4700 0.1750 0.8100 ;
      RECT 0.5950 0.4700 0.6950 0.8100 ;
      RECT 1.1150 0.4700 1.2150 0.8100 ;
      RECT 4.5250 0.5700 4.6250 0.9100 ;
      RECT 1.8550 0.4800 4.6250 0.5700 ;
  END
END NAND3_X6M_A12TH

MACRO NAND4B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.7200 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0100 0.3500 1.3850 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2400 0.5600 1.6250 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.4500 1.1000 1.5700 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8950 1.2400 1.2800 1.3500 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7050 1.5500 1.7000 ;
        RECT 0.6250 1.7000 1.5500 1.8000 ;
        RECT 1.1950 0.6050 1.5500 0.7050 ;
        RECT 0.6250 1.8000 0.7250 1.9800 ;
        RECT 1.1500 1.8000 1.2400 1.9800 ;
        RECT 1.1950 0.5000 1.2950 0.6050 ;
    END
    ANTENNADIFFAREA 0.139375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8500 1.8900 1.0200 2.0800 ;
        RECT 1.3700 1.8900 1.5400 2.0800 ;
        RECT 0.3550 1.7900 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 0.8100 1.3050 0.9000 ;
      RECT 0.0500 1.8700 0.2250 1.9600 ;
      RECT 0.0500 0.9000 0.1400 1.8700 ;
      RECT 0.0500 0.6850 0.1400 0.8100 ;
      RECT 0.0500 0.5950 0.2250 0.6850 ;
  END
END NAND4B_X0P5M_A12TH

MACRO NAND2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1500 0.1600 1.5350 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9950 0.5600 1.3800 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6100 1.7200 0.7100 2.0800 ;
        RECT 0.0900 1.6950 0.1900 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.4750 0.7500 0.9050 ;
        RECT 0.6500 0.9050 0.7500 1.5000 ;
        RECT 0.3500 1.5000 0.7500 1.6000 ;
        RECT 0.3500 1.6000 0.4500 1.9350 ;
    END
    ANTENNADIFFAREA 0.25875 ;
  END Y
END NAND2_X1M_A12TH

MACRO NAND2_X1P4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.7000 ;
        RECT 1.1600 0.3200 1.2600 0.6800 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 1.1500 1.1500 ;
        RECT 1.0600 1.1500 1.1500 1.4200 ;
    END
    ANTENNAGATEAREA 0.1308 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.2500 0.9000 1.3500 ;
    END
    ANTENNAGATEAREA 0.1308 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6450 1.7550 0.7350 2.0800 ;
        RECT 1.1650 1.7550 1.2550 2.0800 ;
        RECT 0.1200 1.6850 0.2200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9000 1.3500 1.5400 ;
        RECT 0.3850 1.5400 1.3500 1.6400 ;
        RECT 0.6400 0.8000 1.3500 0.9000 ;
        RECT 0.3850 1.6400 0.4750 1.9600 ;
        RECT 0.9050 1.6400 0.9950 1.9600 ;
        RECT 0.6400 0.4400 0.7400 0.8000 ;
    END
    ANTENNADIFFAREA 0.327 ;
  END Y
END NAND2_X1P4A_A12TH

MACRO NAND2_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.7500 ;
        RECT 1.1600 0.3200 1.2600 0.7300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 1.1500 1.1500 ;
        RECT 1.0500 1.1500 1.1500 1.4400 ;
    END
    ANTENNAGATEAREA 0.1416 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.2500 0.9100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1416 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6400 1.8400 0.7400 2.0800 ;
        RECT 1.1600 1.8400 1.2600 2.0800 ;
        RECT 0.1200 1.7700 0.2200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.6500 ;
        RECT 0.3450 1.6500 1.3500 1.7500 ;
        RECT 0.6400 0.8500 1.3500 0.9500 ;
        RECT 0.3450 1.7500 0.5150 1.9400 ;
        RECT 0.8650 1.7500 1.0350 1.9400 ;
        RECT 0.6400 0.4450 0.7400 0.8500 ;
    END
    ANTENNADIFFAREA 0.365 ;
  END Y
END NAND2_X1P4B_A12TH

MACRO NAND2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7200 ;
        RECT 1.0250 0.3200 1.1250 0.6900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7550 1.1500 ;
    END
    ANTENNAGATEAREA 0.1182 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.2500 0.9600 1.3500 ;
        RECT 0.8650 1.0100 0.9600 1.2500 ;
    END
    ANTENNAGATEAREA 0.1182 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9000 1.1500 1.4500 ;
        RECT 0.7100 1.4500 1.1500 1.5500 ;
        RECT 0.5250 0.8000 1.1500 0.9000 ;
        RECT 0.7100 1.5500 0.8100 1.9600 ;
        RECT 0.5250 0.4450 0.6250 0.8000 ;
    END
    ANTENNADIFFAREA 0.287725 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4500 1.7500 0.5500 2.0800 ;
        RECT 0.9700 1.7500 1.0700 2.0800 ;
    END
  END VDD
END NAND2_X1P4M_A12TH

MACRO NAND2_X2A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 1.1300 0.3200 1.2300 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 1.0500 1.1500 1.1500 ;
        RECT 1.0500 1.1500 1.1500 1.3000 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.2450 0.9100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.4500 ;
        RECT 0.3500 1.4500 1.3500 1.5500 ;
        RECT 0.6100 0.8500 1.3500 0.9500 ;
        RECT 0.3500 1.5500 0.4500 1.8800 ;
        RECT 0.8700 1.5500 0.9700 1.8800 ;
        RECT 0.6100 0.5200 0.7100 0.8500 ;
    END
    ANTENNADIFFAREA 0.462 ;
  END Y
END NAND2_X2A_A12TH

MACRO NAND2_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1300 0.3200 0.2300 0.6300 ;
        RECT 1.1350 0.3200 1.3050 0.5050 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1300 1.7700 0.2300 2.0800 ;
        RECT 0.6500 1.7700 0.7500 2.0800 ;
        RECT 1.1700 1.7700 1.2700 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 1.1200 1.3500 ;
        RECT 0.2400 1.1500 0.3400 1.2500 ;
        RECT 1.0200 1.0150 1.1200 1.2500 ;
        RECT 0.1300 1.0500 0.3400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1992 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4700 1.0400 0.8900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1992 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7500 1.3500 1.4500 ;
        RECT 0.3900 1.4500 1.3500 1.5500 ;
        RECT 0.6150 0.6500 1.3500 0.7500 ;
        RECT 0.3900 1.5500 0.4900 1.8800 ;
        RECT 0.9100 1.5500 1.0100 1.8800 ;
        RECT 0.6150 0.4600 0.7850 0.6500 ;
    END
    ANTENNADIFFAREA 0.514 ;
  END Y
END NAND2_X2B_A12TH

MACRO NAND2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1300 0.3200 0.2300 0.6300 ;
        RECT 1.1700 0.3200 1.2700 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1300 1.7000 0.2300 2.0800 ;
        RECT 0.6500 1.7000 0.7500 2.0800 ;
        RECT 1.1700 1.7000 1.2700 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1500 1.0500 1.1600 1.1500 ;
        RECT 1.0600 1.1500 1.1600 1.3400 ;
    END
    ANTENNAGATEAREA 0.1668 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.2500 0.9100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1668 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.4500 ;
        RECT 0.3900 1.4500 1.3500 1.5500 ;
        RECT 0.6500 0.8500 1.3500 0.9500 ;
        RECT 0.3900 1.5500 0.4900 1.9400 ;
        RECT 0.9100 1.5500 1.0100 1.9400 ;
        RECT 0.6500 0.5150 0.7500 0.8500 ;
    END
    ANTENNADIFFAREA 0.402 ;
  END Y
END NAND2_X2M_A12TH

MACRO NAND2_X3A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1700 0.3200 0.2700 0.6300 ;
        RECT 1.2100 0.3200 1.3100 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1700 1.7700 0.2700 2.0800 ;
        RECT 0.6900 1.7700 0.7900 2.0800 ;
        RECT 1.2100 1.7700 1.3100 2.0800 ;
        RECT 1.7300 1.7700 1.8300 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.0500 1.5100 1.1500 ;
    END
    ANTENNAGATEAREA 0.2772 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5800 1.2500 1.7500 1.3500 ;
        RECT 1.6500 1.0950 1.7500 1.2500 ;
    END
    ANTENNAGATEAREA 0.2772 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.4500 ;
        RECT 0.4300 1.4500 1.9500 1.5500 ;
        RECT 0.6900 0.8500 1.9500 0.9500 ;
        RECT 0.4300 1.5500 0.5300 1.8800 ;
        RECT 0.9500 1.5500 1.0500 1.8800 ;
        RECT 1.4700 1.5500 1.5700 1.8800 ;
        RECT 0.6900 0.5200 0.7900 0.8500 ;
        RECT 1.7300 0.5200 1.8300 0.8500 ;
    END
    ANTENNADIFFAREA 0.77385 ;
  END Y
END NAND2_X3A_A12TH

MACRO NAND2_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1700 0.3200 0.2700 0.6300 ;
        RECT 1.1750 0.3200 1.3450 0.5050 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1700 1.7700 0.2700 2.0800 ;
        RECT 0.6900 1.7700 0.7900 2.0800 ;
        RECT 1.2100 1.7700 1.3100 2.0800 ;
        RECT 1.7300 1.7700 1.8300 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 0.8500 1.2000 0.9500 ;
        RECT 1.1000 0.9500 1.2000 1.0550 ;
        RECT 0.3000 0.9500 0.4000 1.0500 ;
        RECT 1.1000 1.0550 1.4900 1.1550 ;
        RECT 0.1900 1.0500 0.4000 1.1500 ;
    END
    ANTENNAGATEAREA 0.2988 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8750 1.2500 1.7500 1.3500 ;
        RECT 0.8750 1.1850 0.9750 1.2500 ;
        RECT 1.6500 1.0150 1.7500 1.2500 ;
        RECT 0.5600 1.0850 0.9750 1.1850 ;
    END
    ANTENNAGATEAREA 0.2988 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.7500 1.9500 1.4500 ;
        RECT 0.4300 1.4500 1.9500 1.5500 ;
        RECT 0.6550 0.6500 1.9500 0.7500 ;
        RECT 0.4300 1.5500 0.5300 1.8800 ;
        RECT 0.9500 1.5500 1.0500 1.8800 ;
        RECT 1.4700 1.5500 1.5700 1.8800 ;
        RECT 0.6550 0.4600 0.8250 0.6500 ;
        RECT 1.6950 0.4600 1.8650 0.6500 ;
    END
    ANTENNADIFFAREA 0.84975 ;
  END Y
END NAND2_X3B_A12TH

MACRO NAND2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1700 0.3200 0.2700 0.6300 ;
        RECT 1.2100 0.3200 1.3100 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1700 1.6950 0.2700 2.0800 ;
        RECT 0.6900 1.6950 0.7900 2.0800 ;
        RECT 1.2100 1.6950 1.3100 2.0800 ;
        RECT 1.7300 1.6950 1.8300 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.0500 1.4200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2502 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.2500 1.7500 1.3500 ;
        RECT 1.6500 1.1300 1.7500 1.2500 ;
    END
    ANTENNAGATEAREA 0.2502 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.4500 ;
        RECT 0.4300 1.4500 1.9500 1.5500 ;
        RECT 0.6900 0.8500 1.9500 0.9500 ;
        RECT 0.4300 1.5500 0.5300 1.9350 ;
        RECT 0.9500 1.5500 1.0500 1.9350 ;
        RECT 1.4700 1.5500 1.5700 1.9350 ;
        RECT 0.6900 0.5200 0.7900 0.8500 ;
        RECT 1.7300 0.5200 1.8300 0.8500 ;
    END
    ANTENNADIFFAREA 0.68385 ;
  END Y
END NAND2_X3M_A12TH

MACRO NAND2_X4A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1100 0.3200 0.2100 0.6300 ;
        RECT 1.1500 0.3200 1.2500 0.6300 ;
        RECT 2.1900 0.3200 2.2900 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.1100 1.7700 0.2100 2.0800 ;
        RECT 0.6300 1.7700 0.7300 2.0800 ;
        RECT 1.1500 1.7700 1.2500 2.0800 ;
        RECT 1.6700 1.7700 1.7700 2.0800 ;
        RECT 2.1900 1.7700 2.2900 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0500 2.1400 1.1500 ;
        RECT 2.0400 1.1500 2.1400 1.3050 ;
    END
    ANTENNAGATEAREA 0.3696 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 1.9000 1.3500 ;
    END
    ANTENNAGATEAREA 0.3696 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.4500 ;
        RECT 0.3700 1.4500 2.3500 1.5500 ;
        RECT 0.6300 0.8500 2.3500 0.9500 ;
        RECT 0.3700 1.5500 0.4700 1.8800 ;
        RECT 0.8900 1.5500 0.9900 1.8800 ;
        RECT 1.4100 1.5500 1.5100 1.8800 ;
        RECT 1.9300 1.5500 2.0300 1.8800 ;
        RECT 0.6300 0.5200 0.7300 0.8500 ;
        RECT 1.6700 0.5200 1.7700 0.8500 ;
    END
    ANTENNADIFFAREA 0.924 ;
  END Y
END NAND2_X4A_A12TH

MACRO NAND2_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1100 0.3200 0.2100 0.6300 ;
        RECT 1.1550 0.3200 1.2450 0.5600 ;
        RECT 2.1950 0.3200 2.2850 0.5600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7500 2.3500 1.4550 ;
        RECT 0.3700 1.4550 2.3500 1.5450 ;
        RECT 0.5950 0.6500 2.3500 0.7500 ;
        RECT 0.3700 1.5450 0.4700 1.8850 ;
        RECT 0.8900 1.5450 0.9900 1.8850 ;
        RECT 1.4100 1.5450 1.5100 1.8850 ;
        RECT 1.9300 1.5450 2.0300 1.8850 ;
        RECT 0.5950 0.4600 0.7650 0.6500 ;
        RECT 1.6350 0.4600 1.8050 0.6500 ;
    END
    ANTENNADIFFAREA 1.028 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.1100 1.7700 0.2100 2.0800 ;
        RECT 0.6300 1.7700 0.7300 2.0800 ;
        RECT 1.1500 1.7700 1.2500 2.0800 ;
        RECT 1.6700 1.7700 1.7700 2.0800 ;
        RECT 2.1900 1.7700 2.2900 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.8500 2.1500 0.9500 ;
        RECT 0.2450 0.9500 0.3450 1.0500 ;
        RECT 0.9900 0.9500 1.0900 1.0500 ;
        RECT 2.0400 0.9500 2.1500 1.2250 ;
        RECT 0.1300 1.0500 0.3450 1.1500 ;
        RECT 0.9900 1.0500 1.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.3984 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7600 1.2500 1.6000 1.3500 ;
        RECT 0.7600 1.1500 0.8600 1.2500 ;
        RECT 1.5000 1.1500 1.6000 1.2500 ;
        RECT 0.4700 1.0500 0.8600 1.1500 ;
        RECT 1.5000 1.0500 1.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.3984 ;
  END A
END NAND2_X4B_A12TH

MACRO NAND2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5600 ;
        RECT 1.0900 0.3200 1.1800 0.5600 ;
        RECT 2.0300 0.3200 2.1200 0.6400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0600 0.6500 1.7000 0.7500 ;
        RECT 0.0600 0.7500 0.1500 1.4500 ;
        RECT 0.5600 0.4600 0.7300 0.6500 ;
        RECT 1.5300 0.4100 1.7000 0.6500 ;
        RECT 0.0600 1.4500 1.4700 1.5500 ;
        RECT 0.0600 1.5500 0.9500 1.5600 ;
        RECT 1.3800 1.5500 1.4700 1.8800 ;
        RECT 0.3400 1.5600 0.4300 1.8800 ;
        RECT 0.8600 1.5600 0.9500 1.8800 ;
    END
    ANTENNADIFFAREA 0.806 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7450 0.8500 1.5200 0.9500 ;
        RECT 0.7450 0.9500 0.8550 1.0500 ;
        RECT 1.4100 0.9500 1.5200 1.0500 ;
        RECT 0.4650 1.0500 0.8550 1.1500 ;
        RECT 1.4100 1.0500 1.8200 1.1600 ;
    END
    ANTENNAGATEAREA 0.3342 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 2.0150 1.3500 ;
        RECT 1.9250 1.0700 2.0150 1.2500 ;
        RECT 0.2400 1.0600 0.3300 1.2500 ;
        RECT 0.9500 1.0600 1.3200 1.2500 ;
    END
    ANTENNAGATEAREA 0.3342 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 0.6000 1.7500 0.6900 2.0800 ;
        RECT 1.1200 1.7500 1.2100 2.0800 ;
        RECT 1.6400 1.7500 1.7300 2.0800 ;
    END
  END VDD
END NAND2_X4M_A12TH

MACRO NAND2_X6A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 1.1300 0.3200 1.2300 0.6300 ;
        RECT 2.1700 0.3200 2.2700 0.6300 ;
        RECT 3.2100 0.3200 3.3100 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
        RECT 2.6900 1.7700 2.7900 2.0800 ;
        RECT 3.2100 1.7700 3.3100 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.2500 3.1450 1.3500 ;
        RECT 0.2000 1.1050 0.2900 1.2500 ;
        RECT 3.0350 1.0950 3.1450 1.2500 ;
    END
    ANTENNAGATEAREA 0.5544 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0500 2.9000 1.1500 ;
    END
    ANTENNAGATEAREA 0.5544 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3500 1.4500 3.3500 1.5500 ;
        RECT 0.3500 1.5500 0.4500 1.8800 ;
        RECT 0.8700 1.5500 0.9700 1.8800 ;
        RECT 1.3900 1.5500 1.4900 1.8800 ;
        RECT 1.9100 1.5500 2.0100 1.8800 ;
        RECT 2.4300 1.5500 2.5300 1.8800 ;
        RECT 2.9500 1.5500 3.0500 1.8800 ;
        RECT 3.2500 0.9500 3.3500 1.4500 ;
        RECT 0.6100 0.8500 3.3500 0.9500 ;
        RECT 0.6100 0.5200 0.7100 0.8500 ;
        RECT 1.6500 0.5200 1.7500 0.8500 ;
        RECT 2.6900 0.5200 2.7900 0.8500 ;
    END
    ANTENNADIFFAREA 1.386 ;
  END Y
END NAND2_X6A_A12TH

MACRO NAND2_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 1.0950 0.3200 1.2650 0.5200 ;
        RECT 2.1350 0.3200 2.3050 0.5200 ;
        RECT 3.1850 0.3200 3.3550 0.5200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
        RECT 2.6900 1.7700 2.7900 2.0800 ;
        RECT 3.2100 1.7700 3.3100 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5300 1.0500 2.9100 1.1500 ;
        RECT 2.5300 0.9500 2.6300 1.0500 ;
        RECT 0.7200 0.8500 2.6300 0.9500 ;
        RECT 0.7200 0.9500 0.8200 1.0500 ;
        RECT 1.4900 0.9500 1.5900 1.0500 ;
        RECT 0.4300 1.0500 0.8200 1.1500 ;
        RECT 1.4900 1.0500 1.8600 1.1500 ;
    END
    ANTENNAGATEAREA 0.5976 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5750 0.6500 3.3500 0.7500 ;
        RECT 3.2500 0.7500 3.3500 1.4500 ;
        RECT 0.5750 0.4550 0.7450 0.6500 ;
        RECT 1.6150 0.4550 1.7850 0.6500 ;
        RECT 2.6550 0.4550 2.8250 0.6500 ;
        RECT 0.3500 1.4500 3.3500 1.5500 ;
        RECT 0.3500 1.5500 0.4500 1.8800 ;
        RECT 0.8700 1.5500 0.9700 1.8800 ;
        RECT 1.3900 1.5500 1.4900 1.8800 ;
        RECT 1.9100 1.5500 2.0100 1.8800 ;
        RECT 2.4300 1.5500 2.5300 1.8800 ;
        RECT 2.9500 1.5500 3.0500 1.8800 ;
    END
    ANTENNADIFFAREA 1.542 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.2500 3.1400 1.3500 ;
        RECT 0.2000 1.1500 0.3000 1.2500 ;
        RECT 0.9700 1.1500 1.0700 1.2500 ;
        RECT 2.0100 1.1500 2.1100 1.2500 ;
        RECT 3.0400 1.0150 3.1400 1.2500 ;
        RECT 0.1100 1.0500 0.3000 1.1500 ;
        RECT 0.9700 1.0500 1.3400 1.1500 ;
        RECT 2.0100 1.0500 2.3800 1.1500 ;
    END
    ANTENNAGATEAREA 0.5976 ;
  END B
END NAND2_X6B_A12TH

MACRO NAND2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5700 ;
        RECT 1.1200 0.3200 1.2100 0.5600 ;
        RECT 2.1000 0.3200 2.1900 0.5600 ;
        RECT 3.0300 0.3200 3.1200 0.6000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.6500 2.6900 0.7500 ;
        RECT 0.2500 0.7500 0.3500 0.8500 ;
        RECT 0.5600 0.4100 0.7300 0.6500 ;
        RECT 1.6000 0.4100 1.7700 0.6500 ;
        RECT 2.5200 0.4100 2.6900 0.6500 ;
        RECT 0.0500 0.8500 0.3500 0.9500 ;
        RECT 0.0500 0.9500 0.1500 1.4500 ;
        RECT 0.0500 1.4500 2.5100 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8400 ;
        RECT 0.8600 1.5500 0.9500 1.8400 ;
        RECT 1.3800 1.5500 1.4700 1.8400 ;
        RECT 1.9000 1.5500 1.9900 1.8450 ;
        RECT 2.4200 1.5500 2.5100 1.8450 ;
    END
    ANTENNADIFFAREA 1.207 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0400 2.8200 1.1500 ;
        RECT 0.4650 1.1500 0.8350 1.1600 ;
        RECT 1.5050 1.1500 1.8750 1.1600 ;
    END
    ANTENNAGATEAREA 0.5007 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 3.0600 1.3500 ;
        RECT 0.2500 1.1450 0.3400 1.2500 ;
    END
    ANTENNAGATEAREA 0.5007 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0800 1.8200 0.1700 2.0800 ;
        RECT 0.6000 1.8200 0.6900 2.0800 ;
        RECT 1.1200 1.8200 1.2100 2.0800 ;
        RECT 1.6400 1.8200 1.7300 2.0800 ;
        RECT 2.1600 1.8200 2.2500 2.0800 ;
        RECT 2.6800 1.8200 2.7700 2.0800 ;
    END
  END VDD
END NAND2_X6M_A12TH

MACRO NAND2_X8A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5600 ;
        RECT 1.1200 0.3200 1.2100 0.5600 ;
        RECT 2.1600 0.3200 2.2500 0.5600 ;
        RECT 3.2000 0.3200 3.2900 0.5600 ;
        RECT 4.2300 0.3200 4.3200 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 0.8300 1.1500 ;
        RECT 0.7400 0.9500 0.8300 1.0500 ;
        RECT 0.7400 0.8500 3.6650 0.9500 ;
        RECT 3.5750 0.9500 3.6650 1.0600 ;
        RECT 1.4950 0.9500 2.9150 0.9550 ;
        RECT 3.5750 1.0600 3.9450 1.1500 ;
        RECT 1.4950 0.9550 1.8650 1.1500 ;
        RECT 2.5450 0.9550 2.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.7392 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 4.1650 1.3500 ;
        RECT 0.9750 1.2400 3.4350 1.2500 ;
        RECT 4.0750 1.0700 4.1650 1.2500 ;
        RECT 0.2400 1.0500 0.3300 1.2500 ;
        RECT 0.9750 1.1300 1.3450 1.2400 ;
        RECT 2.0250 1.1100 2.3950 1.2400 ;
        RECT 3.0650 1.1100 3.4350 1.2400 ;
    END
    ANTENNAGATEAREA 0.7392 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 0.0800 1.7600 0.1700 2.0800 ;
        RECT 0.6000 1.7600 0.6900 2.0800 ;
        RECT 1.1200 1.7600 1.2100 2.0800 ;
        RECT 1.6400 1.7600 1.7300 2.0800 ;
        RECT 2.1600 1.7600 2.2500 2.0800 ;
        RECT 2.6800 1.7600 2.7700 2.0800 ;
        RECT 3.2000 1.7600 3.2900 2.0800 ;
        RECT 3.7200 1.7600 3.8100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6500 3.8500 0.7500 ;
        RECT 0.0500 0.7500 0.1500 1.4500 ;
        RECT 0.5600 0.4600 0.7400 0.6500 ;
        RECT 1.6000 0.4100 1.7700 0.6500 ;
        RECT 2.6400 0.4100 2.8100 0.6500 ;
        RECT 3.6800 0.4100 3.8500 0.6500 ;
        RECT 0.0500 1.4500 3.5500 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8800 ;
        RECT 0.8600 1.5500 0.9500 1.8800 ;
        RECT 1.3800 1.5500 1.4700 1.8800 ;
        RECT 1.9000 1.5500 1.9900 1.8800 ;
        RECT 2.4200 1.5500 2.5100 1.8800 ;
        RECT 2.9400 1.5500 3.0300 1.8800 ;
        RECT 3.4600 1.5500 3.5500 1.8800 ;
    END
    ANTENNADIFFAREA 1.848 ;
  END Y
END NAND2_X8A_A12TH

MACRO NAND2_X8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1600 0.3200 0.2600 0.6300 ;
        RECT 1.1650 0.3200 1.3350 0.5200 ;
        RECT 2.2050 0.3200 2.3750 0.5200 ;
        RECT 3.2450 0.3200 3.4150 0.5200 ;
        RECT 4.2850 0.3200 4.4550 0.5200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1600 1.7700 0.2600 2.0800 ;
        RECT 0.6800 1.7700 0.7800 2.0800 ;
        RECT 1.2000 1.7700 1.3000 2.0800 ;
        RECT 1.7200 1.7700 1.8200 2.0800 ;
        RECT 2.2400 1.7700 2.3400 2.0800 ;
        RECT 2.7600 1.7700 2.8600 2.0800 ;
        RECT 3.2800 1.7700 3.3800 2.0800 ;
        RECT 3.8000 1.7700 3.9000 2.0800 ;
        RECT 4.3200 1.7700 4.4200 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6000 1.0500 2.9700 1.1500 ;
        RECT 2.6000 0.9500 2.7000 1.0500 ;
        RECT 0.7900 0.8500 3.7400 0.9500 ;
        RECT 0.7900 0.9500 0.8900 1.0500 ;
        RECT 1.5600 0.9500 1.6600 1.0500 ;
        RECT 3.6400 0.9500 3.7400 1.0500 ;
        RECT 0.5200 1.0500 0.8900 1.1500 ;
        RECT 1.5600 1.0500 1.9300 1.1500 ;
        RECT 3.6400 1.0500 4.0100 1.1500 ;
    END
    ANTENNAGATEAREA 0.7968 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 0.6400 4.5500 0.7600 ;
        RECT 4.4300 0.7600 4.5500 1.4400 ;
        RECT 0.6450 0.4700 0.8150 0.6400 ;
        RECT 1.6850 0.4700 1.8550 0.6400 ;
        RECT 2.7250 0.4700 2.8950 0.6400 ;
        RECT 3.7650 0.4700 3.9350 0.6400 ;
        RECT 0.4200 1.4400 4.5500 1.5600 ;
        RECT 0.4200 1.5600 0.5200 1.8700 ;
        RECT 0.9400 1.5600 1.0400 1.8700 ;
        RECT 1.4600 1.5600 1.5600 1.8700 ;
        RECT 1.9800 1.5600 2.0800 1.8700 ;
        RECT 2.5000 1.5600 2.6000 1.8700 ;
        RECT 3.0200 1.5600 3.1200 1.8700 ;
        RECT 3.5400 1.5600 3.6400 1.8700 ;
        RECT 4.0600 1.5600 4.1600 1.8700 ;
    END
    ANTENNADIFFAREA 2.056 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.2500 4.2650 1.3500 ;
        RECT 0.2900 1.1500 0.3900 1.2500 ;
        RECT 1.0400 1.1500 1.1400 1.2500 ;
        RECT 2.0800 1.1500 2.1800 1.2500 ;
        RECT 3.1200 1.1500 3.2200 1.2500 ;
        RECT 4.1650 1.0150 4.2650 1.2500 ;
        RECT 0.1800 1.0500 0.3900 1.1500 ;
        RECT 1.0400 1.0500 1.4200 1.1500 ;
        RECT 2.0800 1.0500 2.4500 1.1500 ;
        RECT 3.1200 1.0500 3.4900 1.1500 ;
    END
    ANTENNAGATEAREA 0.7968 ;
  END B
END NAND2_X8B_A12TH

MACRO NAND2_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1700 0.3200 0.2700 0.6300 ;
        RECT 1.2100 0.3200 1.3100 0.6300 ;
        RECT 2.2500 0.3200 2.3500 0.6300 ;
        RECT 3.2900 0.3200 3.3900 0.6300 ;
        RECT 4.3300 0.3200 4.4300 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.6900 1.7150 0.7900 2.0800 ;
        RECT 1.2100 1.7150 1.3100 2.0800 ;
        RECT 1.7300 1.7150 1.8300 2.0800 ;
        RECT 2.2500 1.7150 2.3500 2.0800 ;
        RECT 2.7700 1.7150 2.8700 2.0800 ;
        RECT 3.2900 1.7150 3.3900 2.0800 ;
        RECT 3.8100 1.7150 3.9100 2.0800 ;
        RECT 4.3300 1.7150 4.4300 2.0800 ;
        RECT 0.1700 1.6950 0.2700 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.0500 4.0400 1.1500 ;
    END
    ANTENNAGATEAREA 0.6672 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 0.8500 4.5500 0.9500 ;
        RECT 4.4500 0.9500 4.5500 1.4500 ;
        RECT 0.6950 0.5200 0.8050 0.8500 ;
        RECT 1.7300 0.5200 1.8300 0.8500 ;
        RECT 2.7700 0.5200 2.8700 0.8500 ;
        RECT 3.8100 0.5200 3.9100 0.8500 ;
        RECT 0.4300 1.4500 4.5500 1.5500 ;
        RECT 0.4300 1.5500 0.5300 1.9350 ;
        RECT 0.9500 1.5500 1.0500 1.9350 ;
        RECT 1.4700 1.5500 1.5700 1.9350 ;
        RECT 1.9900 1.5500 2.0900 1.9350 ;
        RECT 2.5100 1.5500 2.6100 1.9350 ;
        RECT 3.0300 1.5500 3.1300 1.9350 ;
        RECT 3.5500 1.5500 3.6500 1.9350 ;
        RECT 4.0700 1.5500 4.1700 1.9350 ;
    END
    ANTENNADIFFAREA 1.608 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.2500 4.3500 1.3500 ;
        RECT 4.2500 1.1300 4.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.6672 ;
  END B
END NAND2_X8M_A12TH

MACRO NAND3B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4250 0.3200 0.5250 0.6850 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.0500 0.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.2500 0.7050 1.3500 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6900 1.3500 1.6500 ;
        RECT 0.6900 1.6500 1.3500 1.7500 ;
        RECT 1.1450 0.6000 1.3500 0.6900 ;
        RECT 0.6900 1.7500 0.7800 1.9450 ;
        RECT 1.2100 1.7500 1.3000 1.9450 ;
    END
    ANTENNADIFFAREA 0.15175 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9100 1.8400 1.0800 2.0800 ;
        RECT 0.3600 1.7200 0.4600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5400 1.1450 1.5500 ;
      RECT 0.4800 1.4600 1.1450 1.5400 ;
      RECT 1.0550 0.8750 1.1450 1.4600 ;
      RECT 0.0450 0.7850 1.1450 0.8750 ;
      RECT 0.0950 1.6300 0.1850 1.9450 ;
      RECT 0.0950 1.5500 0.5700 1.6300 ;
  END
END NAND3B_X0P5M_A12TH

MACRO NAND3B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.3900 0.3200 0.5600 0.6650 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9100 1.8400 1.0800 2.0800 ;
        RECT 0.4250 1.7950 0.5250 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6900 1.3500 1.6500 ;
        RECT 0.6900 1.6500 1.3500 1.7500 ;
        RECT 1.1450 0.6000 1.3500 0.6900 ;
        RECT 0.6900 1.7500 0.7800 1.8950 ;
        RECT 1.2100 1.7500 1.3500 1.8950 ;
    END
    ANTENNADIFFAREA 0.215375 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.2500 0.7000 1.3500 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1600 1.3950 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.0500 0.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0519 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.4900 1.4600 1.1450 1.5500 ;
      RECT 1.0550 0.8750 1.1450 1.4600 ;
      RECT 0.0450 0.7850 1.1450 0.8750 ;
      RECT 0.0950 1.6750 0.1850 1.8950 ;
      RECT 0.0950 1.5850 0.5800 1.6750 ;
      RECT 0.4900 1.5500 0.5800 1.5850 ;
  END
END NAND3B_X0P7M_A12TH

MACRO NAND3B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4250 0.3200 0.5250 0.6100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9450 1.8700 1.0450 2.0800 ;
        RECT 0.4300 1.6700 0.5200 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.0100 0.9500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1600 1.3950 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END AN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.2500 0.6750 1.3500 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7150 1.3500 1.6500 ;
        RECT 0.6900 1.6500 1.3500 1.7500 ;
        RECT 1.1700 0.4250 1.3500 0.7150 ;
        RECT 0.6900 1.7500 0.7800 1.8600 ;
        RECT 1.2100 1.7500 1.3500 1.8600 ;
    END
    ANTENNADIFFAREA 0.3035 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2450 1.4600 1.1400 1.5500 ;
      RECT 1.0500 0.9000 1.1400 1.4600 ;
      RECT 0.0450 0.8100 1.1400 0.9000 ;
      RECT 0.0950 1.6200 0.3350 1.7100 ;
      RECT 0.2450 1.5500 0.3350 1.6200 ;
      RECT 0.0950 1.7100 0.1850 1.8300 ;
  END
END NAND3B_X1M_A12TH

MACRO NAND3B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5800 ;
        RECT 1.3550 0.3200 1.4550 0.7050 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.2500 0.9950 1.3500 ;
        RECT 0.9050 1.2400 0.9950 1.2500 ;
        RECT 0.4100 1.1600 0.6000 1.2500 ;
        RECT 0.9050 1.1500 1.1150 1.2400 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 1.4400 1.3100 1.5500 ;
        RECT 1.1000 1.3800 1.3100 1.4400 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0200 1.5500 1.4400 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.6500 1.1800 1.7500 ;
        RECT 0.4900 1.7500 0.6600 1.9550 ;
        RECT 1.0100 1.7500 1.1800 1.9450 ;
        RECT 0.0450 0.7600 0.1350 1.6500 ;
        RECT 0.0450 0.6700 0.8500 0.7600 ;
        RECT 0.6800 0.4500 0.8500 0.6700 ;
    END
    ANTENNADIFFAREA 0.3522 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.7500 1.8600 0.9200 2.0800 ;
        RECT 1.3100 1.7500 1.4000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6300 1.5800 1.7500 1.7900 ;
      RECT 1.6600 0.9000 1.7500 1.5800 ;
      RECT 0.5650 0.8900 1.7500 0.9000 ;
      RECT 0.9450 0.8000 1.7500 0.8900 ;
      RECT 1.6300 0.5550 1.7500 0.8000 ;
      RECT 0.5650 0.9000 1.0550 0.9800 ;
  END
END NAND3B_X1P4M_A12TH

MACRO NAND3B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5600 ;
        RECT 1.5050 0.3200 1.5950 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.2500 1.1500 1.3500 ;
        RECT 0.3000 1.2200 0.5100 1.2500 ;
        RECT 1.0600 1.1800 1.1500 1.2500 ;
        RECT 1.0600 1.0900 1.2700 1.1800 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.4500 1.4900 1.5550 ;
        RECT 1.3900 1.0450 1.4900 1.4500 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6450 1.2400 1.7600 1.6100 ;
    END
    ANTENNAGATEAREA 0.0423 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.6500 1.3750 1.7500 ;
        RECT 0.6850 1.7500 0.8550 1.9600 ;
        RECT 1.2050 1.7500 1.3750 1.9400 ;
        RECT 0.0450 0.7800 0.1350 1.6500 ;
        RECT 0.0450 0.6800 0.8400 0.7800 ;
        RECT 0.7400 0.4100 0.8400 0.6800 ;
    END
    ANTENNADIFFAREA 0.496 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.9450 1.8850 1.1150 2.0800 ;
        RECT 1.5050 1.7600 1.5950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.8200 1.7250 1.9400 1.9350 ;
      RECT 1.8500 0.9550 1.9400 1.7250 ;
      RECT 0.8800 0.8650 1.9400 0.9550 ;
      RECT 1.8300 0.7600 1.9400 0.8650 ;
      RECT 0.8800 0.9550 0.9700 1.0600 ;
      RECT 0.6000 1.0600 0.9700 1.1500 ;
  END
END NAND3B_X2M_A12TH

MACRO NAND3B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.7450 0.3200 0.8350 0.5600 ;
        RECT 2.0650 0.3200 2.1550 0.6300 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8050 0.8500 2.0400 0.9500 ;
        RECT 1.9500 0.9500 2.0400 1.0500 ;
        RECT 0.8050 0.9500 0.9050 1.0450 ;
        RECT 1.9500 1.0500 2.1200 1.1400 ;
        RECT 0.6300 1.0450 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.0500 1.8100 1.1500 ;
        RECT 1.0100 1.1500 1.1150 1.2850 ;
        RECT 1.7100 1.1500 1.8100 1.3600 ;
        RECT 0.4050 1.2850 1.1150 1.3750 ;
    END
    ANTENNAGATEAREA 0.2196 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 1.2500 2.3500 1.3500 ;
        RECT 2.2400 1.1000 2.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.6500 2.0000 1.7150 ;
        RECT 0.0500 1.7150 2.0000 1.7500 ;
        RECT 0.0500 1.7500 0.9600 1.8050 ;
        RECT 1.3100 1.7500 1.4800 1.9500 ;
        RECT 1.8300 1.7500 2.0000 1.9400 ;
        RECT 0.0500 0.7500 0.1500 1.7150 ;
        RECT 0.7900 1.8050 0.9600 1.9500 ;
        RECT 0.0500 0.6500 1.5350 0.7500 ;
        RECT 0.0500 0.5400 0.1700 0.6500 ;
        RECT 1.3650 0.4400 1.5350 0.6500 ;
    END
    ANTENNADIFFAREA 0.6822 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.5300 1.8950 0.7000 2.0800 ;
        RECT 1.0500 1.8800 1.2200 2.0800 ;
        RECT 1.6100 1.8400 1.7000 2.0800 ;
        RECT 2.1300 1.6800 2.2200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2600 1.5600 0.4300 1.6050 ;
      RECT 0.2600 1.4700 2.5500 1.5600 ;
      RECT 2.3900 0.4900 2.4950 0.8200 ;
      RECT 2.3900 0.8200 2.5500 0.9200 ;
      RECT 2.4050 1.5600 2.5050 1.9550 ;
      RECT 2.4600 0.9200 2.5500 1.4700 ;
      RECT 1.3350 1.3350 1.5500 1.5600 ;
  END
END NAND3B_X3M_A12TH

MACRO NAND3B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.1050 0.3200 0.1950 0.6300 ;
        RECT 1.6650 0.3200 1.7550 0.6300 ;
        RECT 3.2250 0.3200 3.3150 0.5700 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 2.9600 1.3500 ;
        RECT 0.4500 1.0700 0.5600 1.2500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4350 0.8500 3.3500 0.9500 ;
        RECT 3.2500 0.9500 3.3500 1.6500 ;
        RECT 2.4350 0.7400 2.5450 0.8500 ;
        RECT 0.0450 1.6500 3.3500 1.7500 ;
        RECT 0.3600 1.7500 0.4600 1.8950 ;
        RECT 0.8800 1.7500 0.9800 1.8950 ;
        RECT 1.4000 1.7500 1.5000 1.8950 ;
        RECT 1.9200 1.7500 2.0200 1.8950 ;
        RECT 2.4400 1.7500 2.5400 1.8950 ;
        RECT 2.9600 1.7500 3.0600 1.8950 ;
        RECT 0.0450 0.9500 0.1500 1.6500 ;
        RECT 0.0450 0.8500 0.9750 0.9500 ;
        RECT 0.8850 0.5200 0.9750 0.8500 ;
    END
    ANTENNADIFFAREA 0.848 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.9100 3.5500 1.3300 ;
    END
    ANTENNAGATEAREA 0.0816 ;
  END AN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.4500 3.1600 1.5500 ;
        RECT 0.2600 1.3500 0.3500 1.4500 ;
        RECT 3.0700 1.3500 3.1600 1.4500 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.1000 1.9250 0.2000 2.0800 ;
        RECT 0.6200 1.9250 0.7200 2.0800 ;
        RECT 1.1400 1.9250 1.2400 2.0800 ;
        RECT 1.6600 1.9250 1.7600 2.0800 ;
        RECT 2.1800 1.9250 2.2800 2.0800 ;
        RECT 2.7000 1.9250 2.8000 2.0800 ;
        RECT 3.2450 1.8600 3.4150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.5600 1.5900 3.6500 1.9300 ;
      RECT 3.5600 1.5000 3.7500 1.5900 ;
      RECT 3.6600 0.7600 3.7500 1.5000 ;
      RECT 2.6800 0.6700 3.7500 0.7600 ;
      RECT 3.5600 0.4300 3.6500 0.6700 ;
      RECT 2.2250 0.5700 2.3150 1.0500 ;
      RECT 0.7700 1.0500 2.3150 1.0550 ;
      RECT 0.7700 1.0550 2.6700 1.1500 ;
      RECT 2.6800 0.5700 2.7700 0.6700 ;
      RECT 2.2250 0.4800 2.7700 0.5700 ;
  END
END NAND3B_X4M_A12TH

MACRO NAND2B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4650 0.3200 0.5550 0.6950 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9450 1.8400 1.1150 2.0800 ;
        RECT 0.4600 1.7500 0.5600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.6750 1.1500 1.6400 ;
        RECT 0.7250 1.6400 1.1500 1.7500 ;
        RECT 0.9150 0.5750 1.1500 0.6750 ;
        RECT 0.7250 1.7500 0.8150 1.8600 ;
    END
    ANTENNADIFFAREA 0.140925 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.2400 0.7100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0417 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1450 1.0300 0.5050 1.1500 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN
  OBS
    LAYER M1 ;
      RECT 0.1300 1.4600 0.9200 1.5500 ;
      RECT 0.8300 0.8750 0.9200 1.4600 ;
      RECT 0.0700 0.7850 0.9200 0.8750 ;
      RECT 0.1300 1.5500 0.2200 1.8550 ;
  END
END NAND2B_X0P5M_A12TH

MACRO NAND2B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4600 0.3200 0.5600 0.6900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9550 1.8650 1.1250 2.0800 ;
        RECT 0.4600 1.7750 0.5600 2.0800 ;
    END
  END VDD

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2250 0.9950 0.3500 1.3700 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5700 1.2100 0.7500 1.3900 ;
        RECT 0.5700 0.9950 0.6600 1.2100 ;
    END
    ANTENNAGATEAREA 0.0591 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.6650 1.1500 1.6600 ;
        RECT 0.6850 1.6600 1.1500 1.7700 ;
        RECT 0.9250 0.5650 1.1500 0.6650 ;
        RECT 0.6850 1.7700 0.8550 1.9900 ;
    END
    ANTENNADIFFAREA 0.187775 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0950 1.4800 0.9300 1.5700 ;
      RECT 0.8400 0.8750 0.9300 1.4800 ;
      RECT 0.0450 0.7850 0.9300 0.8750 ;
      RECT 0.0950 1.5700 0.1850 1.7500 ;
  END
END NAND2B_X0P7M_A12TH

MACRO NAND2B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4650 0.3200 0.5550 0.6300 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.2300 0.3550 1.4050 ;
        RECT 0.0950 1.1200 0.3550 1.2300 ;
    END
    ANTENNAGATEAREA 0.0258 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5700 1.0950 0.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8300 1.1500 1.7050 ;
        RECT 0.6650 1.7050 1.1500 1.8150 ;
        RECT 0.9950 0.7300 1.1500 0.8300 ;
        RECT 0.9950 0.4400 1.0850 0.7300 ;
    END
    ANTENNADIFFAREA 0.26495 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9950 1.9150 1.0850 2.0800 ;
        RECT 0.4650 1.7150 0.5550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1100 1.5050 0.9300 1.5950 ;
      RECT 0.8400 1.0000 0.9300 1.5050 ;
      RECT 0.1100 0.9100 0.9300 1.0000 ;
      RECT 0.1100 1.5950 0.2000 1.7150 ;
      RECT 0.1100 0.7550 0.2000 0.9100 ;
  END
END NAND2B_X1M_A12TH

MACRO NAND2B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3800 0.3200 0.5500 0.7200 ;
        RECT 1.4300 0.3200 1.5200 0.5750 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.2500 1.3500 1.3500 ;
        RECT 1.2500 1.0950 1.3500 1.2500 ;
        RECT 0.4900 1.0700 0.5900 1.2500 ;
    END
    ANTENNAGATEAREA 0.1182 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.4500 ;
        RECT 0.6500 1.4500 1.5500 1.5500 ;
        RECT 0.9100 0.8500 1.5500 0.9500 ;
        RECT 0.6500 1.5500 0.7400 1.8900 ;
        RECT 1.1700 1.5500 1.2600 1.8900 ;
        RECT 0.9100 0.5200 1.0000 0.8500 ;
    END
    ANTENNADIFFAREA 0.285 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3900 1.7100 0.4800 2.0800 ;
        RECT 0.9100 1.7100 1.0000 2.0800 ;
        RECT 1.4300 1.7100 1.5200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.1350 1.1500 ;
      RECT 0.0800 1.5850 0.1700 1.7100 ;
      RECT 0.0800 1.4950 0.3900 1.5850 ;
      RECT 0.3000 0.9000 0.3900 1.4950 ;
      RECT 0.0450 0.8100 0.7900 0.9000 ;
      RECT 0.7000 0.9000 0.7900 1.0600 ;
  END
END NAND2B_X1P4M_A12TH

MACRO NAND2B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3900 0.3200 0.4800 0.6250 ;
        RECT 1.4300 0.3200 1.5200 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3900 1.6700 0.4800 2.0800 ;
        RECT 0.9100 1.6700 1.0000 2.0800 ;
        RECT 1.4300 1.6700 1.5200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9200 1.5500 1.4500 ;
        RECT 0.6500 1.4500 1.5500 1.5500 ;
        RECT 0.9050 0.8200 1.5500 0.9200 ;
        RECT 0.6500 1.5500 0.7400 1.8900 ;
        RECT 1.1700 1.5500 1.2600 1.8900 ;
        RECT 0.9050 0.4900 1.0050 0.8200 ;
    END
    ANTENNADIFFAREA 0.402 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1600 1.4000 ;
    END
    ANTENNAGATEAREA 0.0477 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 1.3500 1.3500 ;
        RECT 0.4500 1.0950 0.5500 1.2500 ;
        RECT 1.2500 1.0950 1.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.1668 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.6550 1.0700 1.1350 1.1600 ;
      RECT 0.0850 1.5850 0.1750 1.9250 ;
      RECT 0.0850 1.4950 0.3450 1.5850 ;
      RECT 0.2550 0.9000 0.3450 1.4950 ;
      RECT 0.0450 0.8100 0.7450 0.9000 ;
      RECT 0.6550 0.9000 0.7450 1.0700 ;
  END
END NAND2B_X2M_A12TH

MACRO NAND2B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6700 ;
        RECT 0.8900 0.3200 0.9800 0.6100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9050 1.9500 1.4500 ;
        RECT 0.6300 1.4500 1.9500 1.5500 ;
        RECT 1.3500 0.8050 2.0200 0.9050 ;
        RECT 0.6300 1.5500 0.7200 1.8950 ;
        RECT 1.1500 1.5500 1.2400 1.8950 ;
        RECT 1.6700 1.5500 1.7600 1.8950 ;
        RECT 1.9300 0.4900 2.0200 0.8050 ;
    END
    ANTENNADIFFAREA 0.68385 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9950 0.3500 1.3850 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6850 1.2500 1.1050 1.3500 ;
    END
    ANTENNAGATEAREA 0.2502 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.8900 1.6850 0.9800 2.0800 ;
        RECT 1.4100 1.6850 1.5000 2.0800 ;
        RECT 1.9300 1.6850 2.0200 2.0800 ;
        RECT 0.3550 1.6650 0.4450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.2900 1.1550 1.7050 1.2550 ;
      RECT 0.4400 1.0500 1.3900 1.1500 ;
      RECT 1.2900 1.1500 1.3900 1.1550 ;
      RECT 0.0950 1.5750 0.1850 1.9150 ;
      RECT 0.0950 0.4700 0.1850 0.7900 ;
      RECT 0.0950 1.4850 0.5300 1.5750 ;
      RECT 0.4400 1.1500 0.5300 1.4850 ;
      RECT 0.4400 0.8800 0.5300 1.0500 ;
      RECT 0.0950 0.7900 0.5300 0.8800 ;
      RECT 1.1500 0.5350 1.8200 0.6250 ;
      RECT 0.6300 0.8550 1.2400 0.9450 ;
      RECT 1.1500 0.6250 1.2400 0.8550 ;
      RECT 0.6300 0.5350 0.7200 0.8550 ;
  END
END NAND2B_X3M_A12TH

MACRO NAND2B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.3850 0.3200 0.4750 0.7150 ;
        RECT 1.3850 0.3200 1.4750 0.6300 ;
        RECT 2.4300 0.3200 2.5200 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.3450 1.7450 0.4350 2.0800 ;
        RECT 0.8650 1.7450 0.9550 2.0800 ;
        RECT 1.3850 1.7450 1.4750 2.0800 ;
        RECT 1.9050 1.7450 1.9950 2.0800 ;
        RECT 2.4250 1.7450 2.5150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9500 2.5500 1.4500 ;
        RECT 0.6050 1.4500 2.5500 1.5500 ;
        RECT 0.8650 0.8500 2.5500 0.9500 ;
        RECT 0.6050 1.5500 0.6950 1.9650 ;
        RECT 1.1250 1.5500 1.2150 1.9650 ;
        RECT 1.6450 1.5500 1.7350 1.9650 ;
        RECT 2.1650 1.5500 2.2550 1.9650 ;
        RECT 0.8650 0.5200 0.9550 0.8500 ;
        RECT 1.9050 0.5200 1.9950 0.8500 ;
    END
    ANTENNADIFFAREA 0.804 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1700 1.3950 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0500 2.3400 1.1500 ;
        RECT 2.2500 1.1500 2.3400 1.3300 ;
    END
    ANTENNAGATEAREA 0.3336 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.2600 1.2600 2.1300 1.3500 ;
      RECT 0.0850 1.5950 0.1750 1.9350 ;
      RECT 0.0850 0.4700 0.1750 0.8100 ;
      RECT 0.0850 1.5050 0.3500 1.5950 ;
      RECT 0.2600 1.3500 0.3500 1.5050 ;
      RECT 0.2600 0.9000 0.3500 1.2600 ;
      RECT 0.0850 0.8100 0.3500 0.9000 ;
  END
END NAND2B_X4M_A12TH

MACRO NAND2B_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.1100 0.3200 0.2000 0.5600 ;
        RECT 1.1200 0.3200 1.2100 0.5600 ;
        RECT 2.1500 0.3200 2.2400 0.5600 ;
        RECT 3.1100 0.3200 3.2000 0.8700 ;
        RECT 3.6300 0.3200 3.7200 0.8900 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2650 1.0700 3.1250 1.1150 ;
        RECT 0.2650 1.1150 0.3550 1.1950 ;
        RECT 0.9750 1.1150 1.3450 1.1800 ;
        RECT 2.0050 1.1150 2.3750 1.1800 ;
        RECT 2.9050 1.1150 3.1250 1.1600 ;
        RECT 0.2650 1.0250 2.9950 1.0700 ;
        RECT 0.2650 0.9850 0.3550 1.0250 ;
    END
    ANTENNAGATEAREA 0.5007 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3950 1.2100 3.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.6500 2.7400 0.7500 ;
        RECT 0.0450 0.7500 0.1500 1.4500 ;
        RECT 0.5900 0.4100 0.7600 0.6500 ;
        RECT 1.6000 0.4100 1.7700 0.6500 ;
        RECT 2.5700 0.4100 2.7400 0.6500 ;
        RECT 0.0450 1.4500 2.5100 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8800 ;
        RECT 0.8600 1.5500 0.9500 1.8800 ;
        RECT 1.3800 1.5500 1.4700 1.8800 ;
        RECT 1.9000 1.5500 1.9900 1.8800 ;
        RECT 2.4200 1.5500 2.5100 1.8800 ;
    END
    ANTENNADIFFAREA 1.207 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.0800 1.8200 0.1700 2.0800 ;
        RECT 0.6000 1.8200 0.6900 2.0800 ;
        RECT 1.1200 1.8200 1.2100 2.0800 ;
        RECT 1.6400 1.8200 1.7300 2.0800 ;
        RECT 2.1600 1.8200 2.2500 2.0800 ;
        RECT 2.6800 1.8200 2.7700 2.0800 ;
        RECT 3.1100 1.7500 3.2000 2.0800 ;
        RECT 3.6300 1.7500 3.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.3700 1.5700 3.4600 1.9100 ;
      RECT 3.2150 1.4800 3.4600 1.5700 ;
      RECT 3.2150 0.9950 3.4600 1.0850 ;
      RECT 3.3700 0.5350 3.4600 0.9950 ;
      RECT 3.2150 1.3600 3.3050 1.4800 ;
      RECT 0.4850 1.2700 3.3050 1.3600 ;
      RECT 3.2150 1.0850 3.3050 1.2700 ;
      RECT 1.5050 1.2050 1.8750 1.2700 ;
      RECT 2.4650 1.2550 2.8350 1.2700 ;
  END
END NAND2B_X6M_A12TH

MACRO NAND2B_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6000 ;
        RECT 1.0000 0.3200 1.0900 0.6000 ;
        RECT 1.9950 0.3200 2.0850 0.6000 ;
        RECT 3.0350 0.3200 3.1250 0.6000 ;
        RECT 4.0150 0.3200 4.1050 0.6000 ;
        RECT 4.5550 0.3200 4.6450 0.6800 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2950 1.0500 4.7350 1.2000 ;
    END
    ANTENNAGATEAREA 0.1836 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1000 1.2500 4.0050 1.3500 ;
        RECT 1.1000 1.2400 1.2500 1.2500 ;
        RECT 1.8500 1.1400 2.2200 1.2500 ;
        RECT 2.8900 1.1400 3.2600 1.2500 ;
        RECT 3.9150 1.1000 4.0050 1.2500 ;
        RECT 0.8350 1.1400 1.2500 1.2400 ;
    END
    ANTENNAGATEAREA 0.6684 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4050 1.4500 3.9050 1.5500 ;
        RECT 1.2150 1.5500 1.3050 1.8800 ;
        RECT 1.7350 1.5500 1.8250 1.8800 ;
        RECT 2.2550 1.5500 2.3450 1.8800 ;
        RECT 2.7750 1.5500 2.8650 1.8800 ;
        RECT 3.2950 1.5500 3.3850 1.8800 ;
        RECT 3.8150 1.5500 3.9050 1.8800 ;
        RECT 0.4050 0.8050 0.5050 1.4500 ;
        RECT 0.4050 0.7050 3.6450 0.8050 ;
        RECT 0.4050 0.7000 0.6300 0.7050 ;
        RECT 1.5350 0.4100 1.6250 0.7050 ;
        RECT 2.5150 0.4100 2.6050 0.7050 ;
        RECT 3.5550 0.4100 3.6450 0.7050 ;
        RECT 0.5400 0.4100 0.6300 0.7000 ;
    END
    ANTENNADIFFAREA 1.612 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.9000 1.7700 0.9900 2.0800 ;
        RECT 1.4750 1.7700 1.5650 2.0800 ;
        RECT 1.9950 1.7700 2.0850 2.0800 ;
        RECT 2.5150 1.7700 2.6050 2.0800 ;
        RECT 3.0350 1.7700 3.1250 2.0800 ;
        RECT 3.5550 1.7700 3.6450 2.0800 ;
        RECT 4.0900 1.7700 4.1800 2.0800 ;
        RECT 4.6100 1.7700 4.7000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.3500 1.3800 4.4400 1.6900 ;
      RECT 4.0950 1.2900 4.4400 1.3800 ;
      RECT 3.7150 0.8650 4.3850 0.9550 ;
      RECT 4.2950 0.5250 4.3850 0.8650 ;
      RECT 4.0950 0.9550 4.1850 1.2900 ;
      RECT 0.6050 1.0500 0.6950 1.1900 ;
      RECT 1.3600 1.0500 1.7300 1.1550 ;
      RECT 2.3800 1.0500 2.7500 1.1550 ;
      RECT 3.3550 1.0500 3.4450 1.0650 ;
      RECT 0.6050 0.9600 3.4450 1.0500 ;
      RECT 3.7150 0.9550 3.8050 1.0650 ;
      RECT 3.3550 1.0650 3.8050 1.1550 ;
  END
END NAND2B_X8M_A12TH

MACRO NAND2XB_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.7300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8350 1.0100 0.9550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0417 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.4150 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9200 1.1500 1.5000 ;
        RECT 0.7300 1.5000 1.1500 1.6100 ;
        RECT 0.9900 0.5100 1.1500 0.9200 ;
        RECT 0.7300 1.6100 0.8200 1.8250 ;
    END
    ANTENNADIFFAREA 0.139 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4650 1.7200 0.5650 2.0800 ;
        RECT 0.9900 1.7200 1.0800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1350 1.5050 0.6250 1.5950 ;
      RECT 0.5350 0.9100 0.6250 1.5050 ;
      RECT 0.0800 0.8200 0.6250 0.9100 ;
      RECT 0.1350 1.5950 0.2250 1.8300 ;
  END
END NAND2XB_X0P5M_A12TH

MACRO NAND2XB_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4500 0.3200 0.6200 0.7350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 1.0050 1.8500 1.1050 2.0800 ;
        RECT 0.4900 1.6600 0.5800 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8650 1.1500 1.6400 ;
        RECT 0.7100 1.6400 1.1500 1.7500 ;
        RECT 1.0100 0.7650 1.1500 0.8650 ;
        RECT 0.7100 1.7500 0.8800 1.9800 ;
        RECT 1.0100 0.4550 1.1000 0.7650 ;
    END
    ANTENNADIFFAREA 0.183375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.0100 0.9600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0591 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END BN
  OBS
    LAYER M1 ;
      RECT 0.1350 1.4800 0.6400 1.5700 ;
      RECT 0.5500 0.9150 0.6400 1.4800 ;
      RECT 0.0750 0.8250 0.6400 0.9150 ;
      RECT 0.1350 1.5700 0.2250 1.8300 ;
  END
END NAND2XB_X0P7M_A12TH

MACRO NAND2XB_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.6300 ;
    END
  END VSS

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0258 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8300 1.0300 0.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9100 1.1500 1.4950 ;
        RECT 0.7300 1.4950 1.1500 1.6050 ;
        RECT 0.9900 0.8100 1.1500 0.9100 ;
        RECT 0.7300 1.6050 0.8200 1.9700 ;
        RECT 0.9900 0.4800 1.0800 0.8100 ;
    END
    ANTENNADIFFAREA 0.278 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4700 1.7500 0.5600 2.0800 ;
        RECT 0.9900 1.7500 1.0800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1150 1.5000 0.6200 1.5900 ;
      RECT 0.5300 0.9200 0.6200 1.5000 ;
      RECT 0.0450 0.8300 0.6200 0.9200 ;
      RECT 0.1150 1.5900 0.2050 1.7700 ;
  END
END NAND2XB_X1M_A12TH

MACRO NAND2XB_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3500 0.3200 0.5200 0.7400 ;
        RECT 1.3250 0.3200 1.4950 0.7400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3900 1.7100 0.4800 2.0800 ;
        RECT 0.9100 1.7100 1.0000 2.0800 ;
        RECT 1.4300 1.7100 1.5200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.4500 ;
        RECT 0.6500 1.4500 1.5500 1.5500 ;
        RECT 0.9100 0.8500 1.5500 0.9500 ;
        RECT 0.6500 1.5500 0.7400 1.9100 ;
        RECT 1.1700 1.5500 1.2600 1.9000 ;
        RECT 0.9100 0.5100 1.0000 0.8500 ;
    END
    ANTENNADIFFAREA 0.285 ;
  END Y

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.0500 1.1350 1.1500 ;
    END
    ANTENNAGATEAREA 0.1182 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4300 1.2500 1.3500 1.3400 ;
      RECT 1.2600 1.0650 1.3500 1.2500 ;
      RECT 0.0800 1.5850 0.1700 1.7100 ;
      RECT 0.0800 0.7000 0.1700 0.8300 ;
      RECT 0.0800 1.4950 0.5200 1.5850 ;
      RECT 0.4300 1.3400 0.5200 1.4950 ;
      RECT 0.4300 0.9200 0.5200 1.2500 ;
      RECT 0.0800 0.8300 0.5200 0.9200 ;
  END
END NAND2XB_X1P4M_A12TH

MACRO NAND2XB_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3900 0.3200 0.4800 0.6300 ;
        RECT 1.4300 0.3200 1.5200 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.0500 1.1350 1.1500 ;
    END
    ANTENNAGATEAREA 0.1668 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0477 ;
  END BN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3900 1.6700 0.4800 2.0800 ;
        RECT 0.9100 1.6650 1.0000 2.0800 ;
        RECT 1.4300 1.6650 1.5200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.4500 ;
        RECT 0.6500 1.4500 1.5500 1.5500 ;
        RECT 0.9100 0.8500 1.5500 0.9500 ;
        RECT 0.6500 1.5500 0.7400 1.9100 ;
        RECT 1.1700 1.5500 1.2600 1.9100 ;
        RECT 0.9100 0.5200 1.0000 0.8500 ;
    END
    ANTENNADIFFAREA 0.402 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.4300 1.2500 1.3500 1.3400 ;
      RECT 1.2600 1.0750 1.3500 1.2500 ;
      RECT 0.0800 1.5700 0.1700 1.9100 ;
      RECT 0.0950 0.7100 0.1850 0.8300 ;
      RECT 0.0800 1.4800 0.5200 1.5700 ;
      RECT 0.4300 1.3400 0.5200 1.4800 ;
      RECT 0.4300 0.9200 0.5200 1.2500 ;
      RECT 0.0950 0.8300 0.5200 0.9200 ;
  END
END NAND2XB_X2M_A12TH

MACRO NAND2XB_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6850 ;
        RECT 0.8900 0.3200 0.9800 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.3550 1.6800 0.4450 2.0800 ;
        RECT 0.8900 1.6550 0.9800 2.0800 ;
        RECT 1.4100 1.6550 1.5000 2.0800 ;
        RECT 1.9300 1.6550 2.0200 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2750 1.0500 1.7050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2502 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9050 1.9500 1.4500 ;
        RECT 0.6300 1.4500 1.9500 1.5500 ;
        RECT 1.3500 0.8050 2.0200 0.9050 ;
        RECT 0.6300 1.5500 0.7200 1.8950 ;
        RECT 1.1500 1.5500 1.2400 1.8950 ;
        RECT 1.6700 1.5500 1.7600 1.8950 ;
        RECT 1.9300 0.4900 2.0200 0.8050 ;
    END
    ANTENNADIFFAREA 0.66075 ;
  END Y

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0300 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END BN
  OBS
    LAYER M1 ;
      RECT 0.4500 1.1550 1.0950 1.2450 ;
      RECT 0.0950 1.5900 0.1850 1.9200 ;
      RECT 0.0950 0.4900 0.1850 0.8300 ;
      RECT 0.0950 1.5000 0.5400 1.5900 ;
      RECT 0.4500 1.2450 0.5400 1.5000 ;
      RECT 0.4500 0.9200 0.5400 1.1550 ;
      RECT 0.0950 0.8300 0.5400 0.9200 ;
      RECT 1.1500 0.4800 1.8250 0.5700 ;
      RECT 0.6300 0.8200 1.2400 0.9100 ;
      RECT 1.1500 0.5700 1.2400 0.8200 ;
      RECT 0.6300 0.4800 0.7200 0.8200 ;
  END
END NAND2XB_X3M_A12TH

MACRO NAND2XB_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.3450 0.3200 0.4350 0.6950 ;
        RECT 1.3850 0.3200 1.4750 0.6300 ;
        RECT 2.4300 0.3200 2.5200 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7300 1.2500 2.1300 1.3500 ;
    END
    ANTENNAGATEAREA 0.3336 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9500 2.5500 1.4500 ;
        RECT 0.6050 1.4500 2.5500 1.5500 ;
        RECT 0.8650 0.8500 2.5500 0.9500 ;
        RECT 0.6050 1.5500 0.6950 1.9650 ;
        RECT 1.1250 1.5500 1.2150 1.9650 ;
        RECT 1.6450 1.5500 1.7350 1.9650 ;
        RECT 2.1650 1.5500 2.2550 1.9650 ;
        RECT 0.8650 0.5200 0.9550 0.8500 ;
        RECT 1.9050 0.5200 1.9950 0.8500 ;
    END
    ANTENNADIFFAREA 0.804 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.8650 1.7650 0.9550 2.0800 ;
        RECT 1.3850 1.7650 1.4750 2.0800 ;
        RECT 1.9050 1.7650 1.9950 2.0800 ;
        RECT 2.4250 1.7650 2.5150 2.0800 ;
        RECT 0.3450 1.7600 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4250 1.0500 2.3600 1.1500 ;
      RECT 2.2700 1.1500 2.3600 1.2750 ;
      RECT 0.0850 1.5700 0.1750 1.9100 ;
      RECT 0.0850 0.4900 0.1750 0.8300 ;
      RECT 0.0850 1.4800 0.5150 1.5700 ;
      RECT 0.4250 1.1500 0.5150 1.4800 ;
      RECT 0.4250 0.9200 0.5150 1.0500 ;
      RECT 0.0850 0.8300 0.5150 0.9200 ;
  END
END NAND2XB_X4M_A12TH

MACRO NAND2XB_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6000 ;
        RECT 1.1200 0.3200 1.2100 0.5600 ;
        RECT 2.1050 0.3200 2.1950 0.5600 ;
        RECT 3.1100 0.3200 3.2000 0.8450 ;
        RECT 3.6300 0.3200 3.7200 0.8200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2650 0.6500 2.7150 0.7500 ;
        RECT 0.2650 0.7500 0.3550 0.9650 ;
        RECT 0.5600 0.4100 0.7300 0.6500 ;
        RECT 1.6000 0.4100 1.7700 0.6500 ;
        RECT 2.5450 0.4100 2.7150 0.6500 ;
        RECT 0.0500 0.9650 0.3550 1.0550 ;
        RECT 0.0500 1.0550 0.1500 1.4500 ;
        RECT 0.0500 1.4500 2.5100 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8400 ;
        RECT 0.8600 1.5500 0.9500 1.8400 ;
        RECT 1.3800 1.5500 1.4700 1.8400 ;
        RECT 1.9000 1.5500 1.9900 1.8450 ;
        RECT 2.4200 1.5500 2.5100 1.8450 ;
    END
    ANTENNADIFFAREA 1.207 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0250 2.8000 1.1250 ;
        RECT 0.4650 1.1250 0.8350 1.1700 ;
        RECT 1.4950 1.1250 1.8650 1.1700 ;
        RECT 2.4050 1.1250 2.8000 1.1500 ;
    END
    ANTENNAGATEAREA 0.5007 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2100 1.2500 3.6300 1.3500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END BN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.0800 1.8200 0.1700 2.0800 ;
        RECT 0.6000 1.8200 0.6900 2.0800 ;
        RECT 1.1200 1.8200 1.2100 2.0800 ;
        RECT 1.6400 1.8200 1.7300 2.0800 ;
        RECT 2.1600 1.8200 2.2500 2.0800 ;
        RECT 2.6800 1.8200 2.7700 2.0800 ;
        RECT 3.1100 1.7650 3.2000 2.0800 ;
        RECT 3.6300 1.7650 3.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.3700 1.5300 3.4600 1.8250 ;
      RECT 2.9300 1.4400 3.4600 1.5300 ;
      RECT 2.9300 0.9950 3.4600 1.0850 ;
      RECT 3.3700 0.6250 3.4600 0.9950 ;
      RECT 0.2600 1.1450 0.3500 1.2600 ;
      RECT 0.9850 1.2500 1.3550 1.2600 ;
      RECT 2.9300 1.3500 3.0300 1.4400 ;
      RECT 0.2600 1.2600 3.0300 1.3500 ;
      RECT 2.9300 1.0850 3.0300 1.2600 ;
  END
END NAND2XB_X6M_A12TH

MACRO NAND2XB_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5600 ;
        RECT 1.0000 0.3200 1.0900 0.5600 ;
        RECT 1.9700 0.3200 2.0600 0.5600 ;
        RECT 3.0100 0.3200 3.1000 0.5600 ;
        RECT 4.0500 0.3200 4.1400 0.6300 ;
        RECT 4.6300 0.3200 4.7200 0.7250 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5450 0.8500 1.4250 0.9500 ;
        RECT 1.3250 0.9500 1.4250 1.0700 ;
        RECT 0.5450 0.9500 0.6350 1.2300 ;
        RECT 1.3250 1.0700 1.6950 1.2000 ;
        RECT 1.5950 0.9550 1.6950 1.0700 ;
        RECT 1.5950 0.8500 3.4750 0.9550 ;
        RECT 3.3850 0.9550 3.4750 1.1100 ;
        RECT 2.3550 0.9550 2.7250 1.2000 ;
        RECT 3.3850 1.1100 3.7550 1.2000 ;
    END
    ANTENNAGATEAREA 0.6684 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2100 1.0500 4.5950 1.2000 ;
    END
    ANTENNAGATEAREA 0.1836 ;
  END BN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6450 3.9200 1.7500 ;
        RECT 1.1800 1.7500 1.2700 1.9900 ;
        RECT 1.7100 1.7500 1.8000 1.9900 ;
        RECT 2.2300 1.7500 2.3200 1.9900 ;
        RECT 2.7500 1.7500 2.8400 1.9900 ;
        RECT 3.2700 1.7500 3.3600 1.9900 ;
        RECT 3.7900 1.7500 3.9200 1.9900 ;
        RECT 0.0500 0.7500 0.1500 1.6450 ;
        RECT 0.0500 0.6500 3.6600 0.7500 ;
        RECT 0.5000 0.4400 0.6700 0.6500 ;
        RECT 1.4300 0.4400 1.6000 0.6500 ;
        RECT 2.4500 0.4400 2.6200 0.6500 ;
        RECT 3.4900 0.4400 3.6600 0.6500 ;
    END
    ANTENNADIFFAREA 1.6203 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.9200 1.8400 1.0100 2.0800 ;
        RECT 1.4500 1.8400 1.5400 2.0800 ;
        RECT 1.9700 1.8400 2.0600 2.0800 ;
        RECT 2.4900 1.8400 2.5800 2.0800 ;
        RECT 3.0100 1.8400 3.1000 2.0800 ;
        RECT 3.5300 1.8400 3.6200 2.0800 ;
        RECT 4.1100 1.7700 4.2000 2.0800 ;
        RECT 4.6300 1.7700 4.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2650 1.2850 0.3550 1.3650 ;
      RECT 0.2650 1.3650 0.9450 1.4550 ;
      RECT 0.8550 1.2300 0.9450 1.3650 ;
      RECT 0.8550 1.1400 1.2250 1.2300 ;
      RECT 1.1250 1.2300 1.2250 1.2900 ;
      RECT 1.1250 1.2900 4.4600 1.3800 ;
      RECT 3.9400 0.8700 4.4200 0.9600 ;
      RECT 3.9400 0.9600 4.0400 1.2900 ;
      RECT 4.3300 0.5800 4.5000 0.8700 ;
      RECT 4.3700 1.3800 4.4600 1.7750 ;
      RECT 1.8250 1.1400 2.1950 1.3800 ;
      RECT 2.8650 1.1400 3.2350 1.3800 ;
  END
END NAND2XB_X8M_A12TH

MACRO NAND2_X0P5A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.7300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7000 0.7500 1.3350 ;
        RECT 0.3500 1.3350 0.7500 1.4350 ;
        RECT 0.5750 0.4100 0.7500 0.7000 ;
        RECT 0.3500 1.4350 0.4500 1.9500 ;
    END
    ANTENNADIFFAREA 0.144375 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.4650 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5550 0.1900 2.0800 ;
        RECT 0.6100 1.5550 0.7100 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.8400 0.5500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END A
END NAND2_X0P5A_A12TH

MACRO NAND2_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.7200 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.4650 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.4200 0.7500 0.7900 ;
        RECT 0.6500 0.7900 0.7500 1.3550 ;
        RECT 0.3500 1.3550 0.7500 1.4450 ;
        RECT 0.3500 1.4450 0.4500 1.9600 ;
    END
    ANTENNADIFFAREA 0.160125 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5850 0.1900 2.0800 ;
        RECT 0.6100 1.5650 0.7100 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.8750 0.5500 1.2600 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END A
END NAND2_X0P5B_A12TH

MACRO NAND2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.7200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7550 0.7500 1.5000 ;
        RECT 0.3500 1.5000 0.7500 1.6000 ;
        RECT 0.5750 0.4250 0.7500 0.7550 ;
        RECT 0.3500 1.6000 0.4500 1.8300 ;
    END
    ANTENNADIFFAREA 0.129375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9950 0.5600 1.3800 ;
    END
    ANTENNAGATEAREA 0.0417 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.7200 0.1900 2.0800 ;
        RECT 0.6100 1.7200 0.7100 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5200 ;
    END
    ANTENNAGATEAREA 0.0417 ;
  END B
END NAND2_X0P5M_A12TH

MACRO NAND2_X0P7A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8350 0.7500 1.5000 ;
        RECT 0.3500 1.5000 0.7500 1.6000 ;
        RECT 0.6150 0.4400 0.7500 0.8350 ;
        RECT 0.3500 1.6000 0.4500 1.9600 ;
    END
    ANTENNADIFFAREA 0.204375 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1850 0.1600 1.5900 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6100 1.7200 0.7100 2.0800 ;
        RECT 0.0900 1.7100 0.1900 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9900 0.5500 1.3750 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END A
END NAND2_X0P7A_A12TH

MACRO NAND2_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7150 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8450 0.7500 1.5000 ;
        RECT 0.3500 1.5000 0.7500 1.6000 ;
        RECT 0.6150 0.4400 0.7500 0.8450 ;
        RECT 0.3500 1.6000 0.4500 1.9350 ;
    END
    ANTENNADIFFAREA 0.222625 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6100 1.6950 0.7100 2.0800 ;
        RECT 0.0900 1.6800 0.1900 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9600 0.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END A
END NAND2_X0P7B_A12TH

MACRO NAND2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7150 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8500 0.7500 1.5000 ;
        RECT 0.3500 1.5000 0.7500 1.6000 ;
        RECT 0.6150 0.4400 0.7500 0.8500 ;
        RECT 0.3500 1.6000 0.4500 1.9900 ;
    END
    ANTENNADIFFAREA 0.183375 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.0591 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6100 1.7000 0.7100 2.0800 ;
        RECT 0.0900 1.6800 0.1900 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9900 0.5500 1.3750 ;
    END
    ANTENNAGATEAREA 0.0591 ;
  END A
END NAND2_X0P7M_A12TH

MACRO NAND2_X1A_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.4850 ;
    END
    ANTENNAGATEAREA 0.0924 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0100 0.5550 1.3950 ;
    END
    ANTENNAGATEAREA 0.0924 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8950 0.7500 1.5150 ;
        RECT 0.3500 1.5150 0.7500 1.6150 ;
        RECT 0.6150 0.4850 0.7500 0.8950 ;
        RECT 0.3500 1.6150 0.4500 1.9450 ;
    END
    ANTENNADIFFAREA 0.28875 ;
  END Y
END NAND2_X1A_A12TH

MACRO NAND2_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6450 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1900 0.1550 1.4100 ;
        RECT 0.0500 1.0800 0.2750 1.1900 ;
    END
    ANTENNAGATEAREA 0.0996 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9950 0.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0996 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.7650 0.1900 2.0800 ;
        RECT 0.6100 1.7650 0.7100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.4600 0.7500 0.8900 ;
        RECT 0.6500 0.8900 0.7500 1.5000 ;
        RECT 0.3500 1.5000 0.7500 1.6000 ;
        RECT 0.3500 1.6000 0.4500 1.9300 ;
    END
    ANTENNADIFFAREA 0.31325 ;
  END Y
END NAND2_X1B_A12TH

MACRO MXIT2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 1.8050 0.3200 1.9050 0.8000 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1400 0.5850 1.4950 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9050 0.3550 1.2200 ;
        RECT 0.2500 0.8050 0.5500 0.9050 ;
        RECT 0.4500 0.5800 0.5500 0.8050 ;
        RECT 0.4500 0.4800 0.9950 0.5800 ;
        RECT 0.8950 0.5800 0.9950 1.0600 ;
        RECT 0.8950 1.0600 1.2150 1.1600 ;
        RECT 1.1250 1.1600 1.2150 1.6150 ;
    END
    ANTENNAGATEAREA 0.1089 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1200 1.8500 1.4300 1.9500 ;
        RECT 1.3300 0.9500 1.4300 1.8500 ;
        RECT 1.1300 0.8500 1.4300 0.9500 ;
        RECT 1.1300 0.4500 1.2200 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1800 1.9500 1.4200 ;
        RECT 1.7250 1.0800 1.9500 1.1800 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.3550 2.0100 0.5250 2.0800 ;
        RECT 1.8050 1.7400 1.9050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7050 0.6900 0.7950 1.7200 ;
      RECT 0.0600 1.8300 0.9850 1.9200 ;
      RECT 0.8950 1.2700 0.9850 1.8300 ;
      RECT 0.0600 0.6850 0.1500 1.8300 ;
      RECT 0.0600 0.5950 0.2300 0.6850 ;
      RECT 1.5450 0.4400 1.6350 1.9600 ;
  END
END MXIT2_X0P7M_A12TH

MACRO MXIT2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 1.8050 0.3200 1.9050 0.6400 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9900 0.5750 1.3900 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8500 0.3600 1.2200 ;
        RECT 0.2500 0.7500 0.5500 0.8500 ;
        RECT 0.4500 0.5800 0.5500 0.7500 ;
        RECT 0.4500 0.4800 1.3500 0.5800 ;
        RECT 1.2500 0.5800 1.3500 1.2700 ;
        RECT 0.8700 0.5800 0.9600 1.1500 ;
        RECT 1.2500 1.2700 1.4300 1.3700 ;
    END
    ANTENNAGATEAREA 0.1482 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.6900 1.1500 1.9300 ;
    END
    ANTENNADIFFAREA 0.45045 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1550 1.9500 1.3900 ;
        RECT 1.7200 1.0550 1.9500 1.1550 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.8050 1.7650 1.9050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6900 0.6900 0.7800 1.6950 ;
      RECT 0.0450 1.8300 0.9600 1.9200 ;
      RECT 0.8700 1.2650 0.9600 1.8300 ;
      RECT 0.0450 1.6200 0.2150 1.8300 ;
      RECT 0.0450 0.5650 0.1350 1.6200 ;
      RECT 0.0450 0.4750 0.2350 0.5650 ;
      RECT 1.5300 0.4700 1.6200 1.9050 ;
  END
END MXIT2_X1M_A12TH

MACRO MXIT2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1600 0.3200 0.2500 0.7050 ;
        RECT 0.6200 0.3200 0.8300 0.3900 ;
        RECT 1.1650 0.3200 1.3750 0.3900 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.0500 0.4650 1.1500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 0.8500 2.3900 0.9500 ;
        RECT 2.2900 0.9500 2.3900 1.0350 ;
        RECT 2.2900 1.0350 2.5450 1.1350 ;
    END
    ANTENNAGATEAREA 0.2022 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7550 0.8500 1.1750 1.0050 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7800 1.4500 3.1500 1.5500 ;
        RECT 2.7800 1.5500 2.8700 1.6400 ;
        RECT 3.0500 0.9200 3.1500 1.4500 ;
        RECT 1.7000 1.6400 2.8700 1.7300 ;
        RECT 3.0300 0.8150 3.1500 0.9200 ;
        RECT 1.7000 1.5900 1.8700 1.6400 ;
        RECT 3.0300 0.5700 3.1200 0.8150 ;
        RECT 1.9300 0.4800 3.1200 0.5700 ;
        RECT 2.5100 0.5700 2.6000 0.8050 ;
        RECT 2.5100 0.4350 2.6000 0.4800 ;
        RECT 3.0300 0.4200 3.1200 0.4800 ;
    END
    ANTENNADIFFAREA 0.5388 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.6800 1.7350 0.7700 2.0800 ;
        RECT 1.2000 1.7350 1.2900 2.0800 ;
        RECT 0.1600 1.4950 0.2500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.5000 1.0500 2.0350 1.1400 ;
      RECT 1.5000 0.6600 1.5900 1.0500 ;
      RECT 1.7250 0.6650 2.4000 0.7550 ;
      RECT 1.1400 1.4100 2.1500 1.5000 ;
      RECT 1.9600 1.5000 2.1500 1.5500 ;
      RECT 0.4200 1.5550 1.2300 1.6450 ;
      RECT 1.1400 1.5000 1.2300 1.5550 ;
      RECT 0.6200 0.4800 1.8150 0.5700 ;
      RECT 1.7250 0.5700 1.8150 0.6650 ;
      RECT 0.4200 1.6450 0.5100 1.9250 ;
      RECT 0.4200 1.5250 0.6450 1.5550 ;
      RECT 0.5550 0.7800 0.6450 1.5250 ;
      RECT 0.4200 0.7600 0.6450 0.7800 ;
      RECT 0.4200 0.4100 0.5100 0.6700 ;
      RECT 0.4200 0.6700 0.7100 0.7600 ;
      RECT 0.6200 0.5700 0.7100 0.6700 ;
      RECT 0.9400 1.2300 2.7800 1.3200 ;
      RECT 2.6900 0.7650 2.7800 1.2300 ;
      RECT 2.6900 0.6600 2.9200 0.7650 ;
      RECT 0.9400 1.3200 1.0300 1.4650 ;
      RECT 1.3000 0.7600 1.3900 1.2300 ;
      RECT 0.8800 0.6700 1.3900 0.7600 ;
      RECT 0.8800 0.6600 1.0900 0.6700 ;
      RECT 2.5200 1.3200 2.6100 1.5100 ;
      RECT 1.4600 1.8600 3.0550 1.9200 ;
      RECT 2.8450 1.9200 3.0550 1.9500 ;
      RECT 1.4600 1.8300 2.9350 1.8600 ;
      RECT 1.5900 1.9200 1.6800 1.9900 ;
      RECT 1.4600 1.8200 1.6800 1.8300 ;
      RECT 1.4600 1.5900 1.5500 1.8200 ;
  END
END MXIT2_X1P4M_A12TH

MACRO MXIT2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.1000 0.3200 0.1900 0.6850 ;
        RECT 0.6200 0.3200 0.7100 0.4500 ;
        RECT 1.1650 0.3200 1.2550 0.4100 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.0500 0.4650 1.1500 ;
    END
    ANTENNAGATEAREA 0.195 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7850 1.1100 1.1550 1.3500 ;
    END
    ANTENNAGATEAREA 0.195 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3000 1.0750 2.7900 1.1500 ;
        RECT 2.7000 1.1500 2.7900 1.1750 ;
        RECT 2.2000 1.0500 2.7900 1.0750 ;
        RECT 2.7000 1.1750 2.9600 1.2750 ;
        RECT 2.2000 0.9850 2.3900 1.0500 ;
    END
    ANTENNAGATEAREA 0.282 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.5800 3.3500 1.5500 ;
        RECT 3.1950 1.5500 3.3500 1.7900 ;
        RECT 2.8650 0.5700 3.3500 0.5800 ;
        RECT 3.1950 1.7900 3.2850 1.8300 ;
        RECT 2.8650 0.5800 2.9550 0.7800 ;
        RECT 1.8250 0.4800 3.3500 0.5700 ;
        RECT 2.1150 1.8300 3.2850 1.9200 ;
        RECT 1.8250 0.5700 1.9150 0.6900 ;
        RECT 2.3450 0.5700 2.4350 0.8500 ;
        RECT 2.8650 0.4100 2.9550 0.4800 ;
    END
    ANTENNADIFFAREA 0.7722 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.2000 2.0100 1.2900 2.0800 ;
        RECT 0.1600 1.7700 0.2500 2.0800 ;
        RECT 0.6800 1.7700 0.7700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6150 1.6500 1.8250 1.7400 ;
      RECT 1.6150 1.3650 1.7050 1.6500 ;
      RECT 1.4250 1.2750 1.9100 1.3650 ;
      RECT 1.4250 1.3650 1.5150 1.6700 ;
      RECT 1.8200 1.1550 1.9100 1.2750 ;
      RECT 1.4250 0.7400 1.5150 1.2750 ;
      RECT 2.0000 1.4100 2.5550 1.5000 ;
      RECT 0.5550 0.5400 1.7150 0.6300 ;
      RECT 1.6250 0.6300 1.7150 0.8050 ;
      RECT 2.0000 0.8950 2.0900 1.4100 ;
      RECT 1.6250 0.8050 2.1750 0.8950 ;
      RECT 2.0850 0.6700 2.1750 0.8050 ;
      RECT 0.4200 1.5300 0.5100 1.8700 ;
      RECT 0.4200 1.4400 0.6450 1.5300 ;
      RECT 0.5550 0.9400 0.6450 1.4400 ;
      RECT 0.3600 0.8500 0.6450 0.9400 ;
      RECT 0.5550 0.6300 0.6450 0.8500 ;
      RECT 0.3600 0.5500 0.4500 0.8500 ;
      RECT 1.9350 1.5900 3.0250 1.6800 ;
      RECT 2.9350 1.4550 3.0250 1.5900 ;
      RECT 2.9350 1.3650 3.1600 1.4550 ;
      RECT 3.0700 0.9600 3.1600 1.3650 ;
      RECT 2.6050 0.8700 3.1600 0.9600 ;
      RECT 1.2450 1.8300 2.0250 1.9200 ;
      RECT 1.9350 1.6800 2.0250 1.8300 ;
      RECT 1.2450 1.5900 1.3350 1.8300 ;
      RECT 0.9400 1.5000 1.3350 1.5900 ;
      RECT 0.9400 1.5900 1.0300 1.9300 ;
      RECT 1.2450 1.0150 1.3350 1.5000 ;
      RECT 0.8800 0.9250 1.3350 1.0150 ;
      RECT 0.8800 0.7400 0.9700 0.9250 ;
      RECT 2.6050 0.6950 2.6950 0.8700 ;
  END
END MXIT2_X2M_A12TH

MACRO MXIT2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.1150 0.3200 0.2150 0.6300 ;
        RECT 0.6350 0.3200 0.7350 0.6300 ;
        RECT 1.1550 0.3200 1.2550 0.6300 ;
        RECT 3.3300 0.3200 3.5000 0.3900 ;
        RECT 3.8500 0.3200 4.0200 0.3900 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2300 1.0500 3.6800 1.1500 ;
    END
    ANTENNAGATEAREA 0.2925 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.5800 4.1500 1.8200 ;
        RECT 1.6200 1.8200 4.1500 1.9200 ;
        RECT 1.6200 0.4800 4.1500 0.5800 ;
    END
    ANTENNADIFFAREA 1.0439 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8650 1.0500 1.2850 1.1500 ;
    END
    ANTENNAGATEAREA 0.2925 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.2500 1.9600 1.3500 ;
        RECT 0.5600 1.0200 0.6500 1.2500 ;
    END
    ANTENNAGATEAREA 0.4134 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 3.3300 2.0300 3.5000 2.0800 ;
        RECT 3.8500 2.0300 4.0200 2.0800 ;
        RECT 1.1550 1.8200 1.2550 2.0800 ;
        RECT 0.1150 1.7700 0.2150 2.0800 ;
        RECT 0.6350 1.7700 0.7350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8600 1.6250 2.4000 1.7150 ;
      RECT 2.3100 1.5400 2.4000 1.6250 ;
      RECT 2.3100 1.4500 3.0700 1.5400 ;
      RECT 2.9800 1.1200 3.0700 1.4500 ;
      RECT 2.3100 1.0300 3.0700 1.1200 ;
      RECT 2.3100 0.8200 2.4000 1.0300 ;
      RECT 0.8400 0.7300 2.4000 0.8200 ;
      RECT 0.8600 1.7150 1.0300 1.9700 ;
      RECT 2.5300 1.6300 3.7200 1.7200 ;
      RECT 3.6300 1.3800 3.7200 1.6300 ;
      RECT 3.6300 1.2900 3.9400 1.3800 ;
      RECT 3.8500 0.7900 3.9400 1.2900 ;
      RECT 2.5300 0.7000 3.9400 0.7900 ;
      RECT 0.3800 1.4450 2.1600 1.5350 ;
      RECT 2.0700 1.3500 2.1600 1.4450 ;
      RECT 2.0700 1.2600 2.8650 1.3500 ;
      RECT 2.0700 1.1050 2.1600 1.2600 ;
      RECT 1.6500 1.0150 2.1600 1.1050 ;
      RECT 0.3800 1.5350 0.4700 1.8600 ;
      RECT 0.3800 0.4900 0.4700 1.4450 ;
  END
END MXIT2_X3M_A12TH

MACRO MXIT2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.3750 0.3200 0.4750 0.6300 ;
        RECT 0.9150 0.3200 1.0150 0.6300 ;
        RECT 1.4350 0.3200 1.5350 0.6300 ;
        RECT 1.9700 0.3200 2.0700 0.6300 ;
        RECT 4.7100 0.3200 4.8800 0.3900 ;
        RECT 5.2300 0.3200 5.4000 0.3900 ;
        RECT 5.7500 0.3200 5.9200 0.3900 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9200 1.0500 5.3900 1.1500 ;
    END
    ANTENNAGATEAREA 0.39 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.5800 5.9500 1.8200 ;
        RECT 2.1900 1.8200 5.9500 1.9200 ;
        RECT 2.1900 0.4800 5.9500 0.5800 ;
    END
    ANTENNADIFFAREA 1.5587 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1450 1.0500 1.7950 1.1500 ;
    END
    ANTENNAGATEAREA 0.39 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6650 1.2500 3.0500 1.3500 ;
        RECT 0.6650 1.1600 0.7550 1.2500 ;
        RECT 0.3350 1.0700 0.7550 1.1600 ;
    END
    ANTENNAGATEAREA 0.5475 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 4.7100 2.0100 4.8800 2.0800 ;
        RECT 5.2300 2.0100 5.4000 2.0800 ;
        RECT 5.7500 2.0100 5.9200 2.0800 ;
        RECT 1.4400 1.8100 1.5300 2.0800 ;
        RECT 1.9600 1.8100 2.0500 2.0800 ;
        RECT 0.3750 1.7700 0.4750 2.0800 ;
        RECT 0.9150 1.7700 1.0150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1200 1.4450 3.2500 1.5350 ;
      RECT 3.1600 1.3500 3.2500 1.4450 ;
      RECT 3.1600 1.2600 4.2950 1.3500 ;
      RECT 3.1600 1.1050 3.2500 1.2600 ;
      RECT 2.4700 1.0150 3.2500 1.1050 ;
      RECT 0.1200 1.5350 0.2100 1.9700 ;
      RECT 0.1200 0.8950 0.2100 1.4450 ;
      RECT 0.1200 0.4550 0.2100 0.8050 ;
      RECT 0.6500 1.5350 0.7400 1.9500 ;
      RECT 0.1200 0.8050 0.7400 0.8950 ;
      RECT 0.6500 0.4550 0.7400 0.8050 ;
      RECT 1.1400 1.6250 3.4750 1.7150 ;
      RECT 3.3850 1.5400 3.4750 1.6250 ;
      RECT 3.3850 1.4500 4.4950 1.5400 ;
      RECT 4.4050 1.1200 4.4950 1.4500 ;
      RECT 3.4000 1.0300 4.4950 1.1200 ;
      RECT 3.4000 0.8300 3.4900 1.0300 ;
      RECT 1.1750 0.7400 3.4900 0.8300 ;
      RECT 1.1400 1.7150 1.3100 1.9700 ;
      RECT 1.1750 0.4400 1.2750 0.7400 ;
      RECT 1.7000 1.7150 1.7900 1.9900 ;
      RECT 1.6950 0.4400 1.7950 0.7400 ;
      RECT 3.6200 1.6300 5.6200 1.7200 ;
      RECT 5.0100 1.3000 5.1000 1.6300 ;
      RECT 5.5300 0.7800 5.6200 1.6300 ;
      RECT 3.6200 0.6900 5.7000 0.7800 ;
  END
END MXIT2_X4M_A12TH

MACRO MXIT4_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.4250 0.3200 0.5150 0.3950 ;
        RECT 1.7650 0.3200 1.8550 0.3950 ;
        RECT 2.2300 0.3200 2.3200 0.7600 ;
        RECT 3.6750 0.3200 3.7650 0.4600 ;
        RECT 5.1000 0.3200 5.1900 0.4600 ;
    END
  END VSS

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0100 2.1500 1.2050 ;
        RECT 2.0500 0.5750 2.1400 1.0100 ;
        RECT 1.1850 0.4850 2.1400 0.5750 ;
        RECT 1.1850 0.5750 1.2750 0.8450 ;
        RECT 0.8500 0.8450 1.3500 0.9350 ;
        RECT 1.2600 0.9350 1.3500 1.0500 ;
        RECT 0.8500 0.9350 0.9400 1.0550 ;
        RECT 1.2600 1.0500 1.4700 1.1400 ;
    END
    ANTENNAGATEAREA 0.0537 ;
  END S1

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.2050 2.3500 1.4150 ;
        RECT 2.2500 1.1150 2.4700 1.2050 ;
        RECT 2.3800 0.9950 2.4700 1.1150 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.7650 3.5550 1.2750 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8250 0.9950 4.0250 1.2050 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0350 0.9950 5.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.4100 5.3400 1.5000 ;
        RECT 5.0500 1.5000 5.1500 1.7600 ;
        RECT 5.2500 1.2800 5.3400 1.4100 ;
        RECT 4.6750 1.7600 5.1500 1.7900 ;
        RECT 3.4000 1.7900 5.1500 1.8500 ;
        RECT 4.6750 1.2150 4.7650 1.7600 ;
        RECT 3.4000 1.8500 4.7650 1.8800 ;
        RECT 3.4000 1.8800 3.4900 1.9000 ;
        RECT 3.3000 1.9000 3.4900 1.9900 ;
    END
    ANTENNAGATEAREA 0.1182 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 0.8100 0.3500 0.9900 ;
        RECT 0.0800 0.9900 0.1700 1.8550 ;
        RECT 0.0800 0.6900 0.1750 0.8100 ;
        RECT 0.0850 0.4100 0.1750 0.6900 ;
    END
    ANTENNADIFFAREA 0.13365 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 2.2300 2.0200 2.3200 2.0800 ;
        RECT 1.7750 2.0100 1.8650 2.0800 ;
        RECT 3.7650 1.9700 3.8550 2.0800 ;
        RECT 5.1500 1.9400 5.2400 2.0800 ;
        RECT 0.4050 1.8200 0.4950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6200 0.6650 0.8950 0.7550 ;
      RECT 0.6200 1.4400 0.8200 1.5300 ;
      RECT 0.6200 0.7550 0.7100 1.4400 ;
      RECT 0.4400 0.5750 0.5300 1.1350 ;
      RECT 0.4400 1.3450 0.5300 1.6400 ;
      RECT 0.4400 0.4850 1.0950 0.5750 ;
      RECT 0.4400 1.6400 1.1150 1.7300 ;
      RECT 1.0050 0.5750 1.0950 0.6950 ;
      RECT 1.0250 1.5400 1.1150 1.6400 ;
      RECT 0.2600 1.1350 0.5300 1.3450 ;
      RECT 1.4550 1.3700 1.5450 1.5400 ;
      RECT 1.4550 1.2800 1.6500 1.3700 ;
      RECT 1.5600 0.7550 1.6500 1.2800 ;
      RECT 1.3850 0.6650 1.6500 0.7550 ;
      RECT 1.2250 1.6500 1.7250 1.7400 ;
      RECT 1.6350 1.5500 1.7250 1.6500 ;
      RECT 1.2250 1.4500 1.3150 1.6500 ;
      RECT 1.6350 1.4600 1.9900 1.5500 ;
      RECT 1.1000 1.3600 1.3150 1.4500 ;
      RECT 1.8700 1.3550 1.9900 1.4600 ;
      RECT 1.8700 0.7150 1.9600 1.3550 ;
      RECT 1.1000 1.3200 1.1900 1.3600 ;
      RECT 0.8000 1.2300 1.1900 1.3200 ;
      RECT 2.5100 1.4200 2.6000 1.5500 ;
      RECT 2.5100 1.3300 2.6500 1.4200 ;
      RECT 2.5600 0.7300 2.6500 1.3300 ;
      RECT 1.8150 1.6400 3.0100 1.7300 ;
      RECT 2.9200 0.7500 3.0100 1.6400 ;
      RECT 0.6300 1.9200 0.8400 1.9900 ;
      RECT 0.6300 1.9000 1.9050 1.9200 ;
      RECT 0.7500 1.8300 1.9050 1.9000 ;
      RECT 1.8150 1.7300 1.9050 1.8300 ;
      RECT 3.2700 0.7500 3.3600 1.5200 ;
      RECT 4.0850 1.4200 4.1750 1.5200 ;
      RECT 4.0850 1.3300 4.2050 1.4200 ;
      RECT 4.1150 0.7500 4.2050 1.3300 ;
      RECT 3.1000 1.6100 4.5850 1.7000 ;
      RECT 4.4950 0.7300 4.5850 1.6100 ;
      RECT 1.9950 1.8400 3.1900 1.9200 ;
      RECT 2.0950 1.8300 3.1900 1.8400 ;
      RECT 3.1000 1.7000 3.1900 1.8300 ;
      RECT 1.9950 1.9200 2.1850 1.9300 ;
      RECT 4.8550 0.9400 4.9450 1.6500 ;
      RECT 4.7550 0.8500 4.9450 0.9400 ;
      RECT 4.7550 0.7300 4.8450 0.8500 ;
      RECT 2.7400 0.6400 2.8300 1.4950 ;
      RECT 2.7400 0.5500 5.5200 0.6400 ;
      RECT 4.2950 0.6400 4.3850 1.2850 ;
      RECT 4.2950 1.2850 4.4050 1.3750 ;
      RECT 4.3150 1.3750 4.4050 1.4950 ;
      RECT 5.4300 1.5850 5.5200 1.9050 ;
      RECT 5.4300 1.4950 5.5500 1.5850 ;
      RECT 5.4300 0.7650 5.5500 0.8550 ;
      RECT 5.4300 0.6400 5.5200 0.7650 ;
      RECT 5.4500 0.8550 5.5500 1.4950 ;
      RECT 2.8650 0.4100 3.0750 0.6400 ;
      RECT 4.5100 0.4100 4.7200 0.6400 ;
  END
END MXIT4_X0P5M_A12TH

MACRO MXIT4_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3950 0.3200 0.5650 0.3850 ;
        RECT 2.0350 0.3200 2.1350 0.6800 ;
        RECT 3.4550 0.3200 3.6250 0.3900 ;
        RECT 3.9800 0.3200 4.1500 0.3900 ;
        RECT 5.3300 0.3200 5.5000 0.5600 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1800 0.5500 1.3900 ;
        RECT 0.4500 0.9900 0.5900 1.1800 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3600 1.2200 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3900 1.1700 3.5600 1.3400 ;
        RECT 3.4500 1.3400 3.5600 1.5500 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9900 1.0500 2.4150 1.1500 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7750 0.8500 2.5350 0.9500 ;
        RECT 1.7750 0.9500 1.8750 1.1800 ;
    END
    ANTENNAGATEAREA 0.1368 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9300 1.0500 5.3000 1.1500 ;
        RECT 5.1800 1.1500 5.3000 1.3000 ;
    END
    ANTENNAGATEAREA 0.0624 ;
  END S1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6300 0.5150 5.7500 1.8250 ;
    END
    ANTENNADIFFAREA 0.1816 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 1.9850 2.0250 2.1550 2.0800 ;
        RECT 3.9750 1.9150 4.1650 2.0800 ;
        RECT 3.4450 1.8800 3.6200 2.0800 ;
        RECT 0.3450 1.6800 0.4350 2.0800 ;
        RECT 5.3650 1.4500 5.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5250 1.8050 1.1000 1.8950 ;
      RECT 0.5250 1.5700 0.6150 1.8050 ;
      RECT 0.0600 1.4800 0.6150 1.5700 ;
      RECT 0.0600 0.4800 1.6450 0.5700 ;
      RECT 0.0600 1.5700 0.1750 1.8800 ;
      RECT 0.0600 0.5700 0.1500 1.4800 ;
      RECT 1.2100 1.8050 1.6500 1.8950 ;
      RECT 1.2100 1.7150 1.3000 1.8050 ;
      RECT 0.7050 1.6250 1.3000 1.7150 ;
      RECT 0.7050 0.7900 0.7950 1.6250 ;
      RECT 0.6650 0.7000 1.0850 0.7900 ;
      RECT 2.3000 1.3300 2.3900 1.5350 ;
      RECT 2.3000 1.2400 2.7350 1.3300 ;
      RECT 2.6450 0.7500 2.7350 1.2400 ;
      RECT 2.3000 0.6600 2.7350 0.7500 ;
      RECT 2.3000 0.5100 2.3900 0.6600 ;
      RECT 2.0550 1.6450 2.5700 1.7350 ;
      RECT 2.0550 1.5350 2.1450 1.6450 ;
      RECT 2.4800 1.5100 2.5700 1.6450 ;
      RECT 1.6200 1.4450 2.1450 1.5350 ;
      RECT 2.4800 1.4200 2.9150 1.5100 ;
      RECT 2.8250 0.8500 2.9150 1.4200 ;
      RECT 1.5300 0.6600 1.8450 0.7500 ;
      RECT 1.7550 0.4850 1.8450 0.6600 ;
      RECT 1.6200 1.3550 1.7100 1.4450 ;
      RECT 1.1550 1.2650 1.7100 1.3550 ;
      RECT 1.1550 1.1450 1.2450 1.2650 ;
      RECT 1.5300 0.7500 1.6200 1.2650 ;
      RECT 3.1850 1.4800 3.3550 1.5700 ;
      RECT 3.1850 0.7700 3.2750 1.4800 ;
      RECT 3.1850 0.6800 3.3750 0.7700 ;
      RECT 2.6050 0.4800 3.6800 0.5700 ;
      RECT 3.5900 0.5700 3.6800 1.0550 ;
      RECT 2.6800 1.6300 3.0950 1.7200 ;
      RECT 3.0050 0.5700 3.0950 1.6300 ;
      RECT 3.2500 1.7000 4.0600 1.7900 ;
      RECT 3.9700 1.0850 4.0600 1.7000 ;
      RECT 1.8550 1.8300 3.3400 1.9200 ;
      RECT 3.2500 1.7900 3.3400 1.8300 ;
      RECT 1.8550 1.7150 1.9450 1.8300 ;
      RECT 1.4100 1.6250 1.9450 1.7150 ;
      RECT 1.4100 1.5350 1.5000 1.6250 ;
      RECT 0.9150 1.4450 1.5000 1.5350 ;
      RECT 0.9150 1.0350 1.0050 1.4450 ;
      RECT 0.9150 0.9450 1.2800 1.0350 ;
      RECT 1.1900 0.7850 1.2800 0.9450 ;
      RECT 1.1900 0.6950 1.3800 0.7850 ;
      RECT 4.3300 0.6600 4.4200 1.5950 ;
      RECT 4.1500 1.7050 4.9800 1.7950 ;
      RECT 4.8100 1.6350 4.9800 1.7050 ;
      RECT 3.7700 0.4800 5.0000 0.5700 ;
      RECT 4.7850 0.5700 5.0000 0.5800 ;
      RECT 4.1500 0.9700 4.2400 1.7050 ;
      RECT 3.7700 0.8800 4.2400 0.9700 ;
      RECT 3.7700 0.9700 3.8600 1.6100 ;
      RECT 3.7700 0.5700 3.8600 0.8800 ;
      RECT 4.8700 1.4550 5.2500 1.5450 ;
      RECT 4.7300 0.8500 5.1900 0.9400 ;
      RECT 4.7300 0.9400 4.8200 1.2400 ;
      RECT 4.8700 1.3300 4.9600 1.4550 ;
      RECT 4.7300 1.2400 4.9600 1.3300 ;
      RECT 4.5300 0.6700 5.5350 0.7600 ;
      RECT 5.4450 0.7600 5.5350 1.2300 ;
      RECT 4.5300 1.4700 4.7400 1.5600 ;
      RECT 4.5300 0.7600 4.6200 1.4700 ;
  END
END MXIT4_X0P7M_A12TH

MACRO MXIT4_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3950 0.3200 0.5650 0.3850 ;
        RECT 2.0350 0.3200 2.1350 0.7400 ;
        RECT 4.0000 0.3200 4.1700 0.3900 ;
        RECT 5.3300 0.3200 5.5000 0.4200 ;
    END
  END VSS

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7750 0.8500 2.5400 0.9500 ;
        RECT 1.7750 0.9500 1.8750 1.1800 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END S0

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9900 1.0500 2.4150 1.1500 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1800 0.5500 1.3900 ;
        RECT 0.4500 0.9900 0.5900 1.1800 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3600 1.2200 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4300 1.1700 3.5500 1.5500 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END C

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8950 1.0500 5.2750 1.1500 ;
        RECT 5.1850 1.1500 5.2750 1.2600 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END S1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6300 0.5250 5.7500 1.7500 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 1.9850 2.0250 2.1550 2.0800 ;
        RECT 5.3700 2.0150 5.4600 2.0800 ;
        RECT 3.4500 1.9150 3.6400 2.0800 ;
        RECT 3.9900 1.9150 4.1800 2.0800 ;
        RECT 0.3450 1.6800 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5250 1.8050 1.1000 1.8950 ;
      RECT 0.5250 1.5700 0.6150 1.8050 ;
      RECT 0.0600 1.4800 0.6150 1.5700 ;
      RECT 0.0600 0.4800 1.6450 0.5700 ;
      RECT 0.0600 1.5700 0.1750 1.8800 ;
      RECT 0.0600 0.5700 0.1500 1.4800 ;
      RECT 1.2100 1.8050 1.6500 1.8950 ;
      RECT 1.2100 1.7150 1.3000 1.8050 ;
      RECT 0.7050 1.6250 1.3000 1.7150 ;
      RECT 0.7050 0.7900 0.7950 1.6250 ;
      RECT 0.7050 0.7000 1.1000 0.7900 ;
      RECT 2.3000 1.3300 2.3900 1.5350 ;
      RECT 2.3000 1.2400 2.7400 1.3300 ;
      RECT 2.6500 0.7500 2.7400 1.2400 ;
      RECT 2.3000 0.6600 2.7400 0.7500 ;
      RECT 2.3000 0.5100 2.3900 0.6600 ;
      RECT 2.0550 1.6450 2.5700 1.7350 ;
      RECT 2.0550 1.5350 2.1450 1.6450 ;
      RECT 2.4800 1.5200 2.5700 1.6450 ;
      RECT 1.6200 1.4450 2.1450 1.5350 ;
      RECT 2.4800 1.4300 2.9200 1.5200 ;
      RECT 2.8300 0.8500 2.9200 1.4300 ;
      RECT 1.5300 0.6600 1.8450 0.7500 ;
      RECT 1.7550 0.4850 1.8450 0.6600 ;
      RECT 1.6200 1.3550 1.7100 1.4450 ;
      RECT 1.1550 1.2650 1.7100 1.3550 ;
      RECT 1.1550 1.1450 1.2450 1.2650 ;
      RECT 1.5300 0.7500 1.6200 1.2650 ;
      RECT 3.1900 0.7750 3.2800 1.6250 ;
      RECT 3.1900 0.6850 3.3800 0.7750 ;
      RECT 2.6050 0.4800 3.6800 0.5700 ;
      RECT 3.5900 0.5700 3.6800 1.0550 ;
      RECT 2.6600 1.6300 3.1000 1.7200 ;
      RECT 3.0100 0.5700 3.1000 1.6300 ;
      RECT 3.2500 1.7350 4.0400 1.8250 ;
      RECT 3.9500 1.0850 4.0400 1.7350 ;
      RECT 1.8550 1.8300 3.3400 1.9200 ;
      RECT 3.2500 1.8250 3.3400 1.8300 ;
      RECT 1.8550 1.7150 1.9450 1.8300 ;
      RECT 1.4100 1.6250 1.9450 1.7150 ;
      RECT 1.4100 1.5350 1.5000 1.6250 ;
      RECT 0.9150 1.4450 1.5000 1.5350 ;
      RECT 0.9150 1.0350 1.0050 1.4450 ;
      RECT 0.9150 0.9450 1.2800 1.0350 ;
      RECT 1.1900 0.7500 1.2800 0.9450 ;
      RECT 1.1900 0.6600 1.3800 0.7500 ;
      RECT 4.3150 0.6600 4.4050 1.6150 ;
      RECT 4.1300 1.7250 4.9850 1.8150 ;
      RECT 3.7700 0.4800 4.9850 0.5700 ;
      RECT 4.1300 0.9750 4.2200 1.7250 ;
      RECT 3.7700 0.8850 4.2200 0.9750 ;
      RECT 3.7700 0.9750 3.8600 1.6250 ;
      RECT 3.7700 0.5700 3.8600 0.8850 ;
      RECT 3.7700 0.4300 3.8600 0.4800 ;
      RECT 4.8150 1.3900 5.2500 1.4800 ;
      RECT 4.6950 0.8700 5.2100 0.9600 ;
      RECT 5.0400 0.8600 5.2100 0.8700 ;
      RECT 4.6950 0.9600 4.7850 1.2400 ;
      RECT 4.8150 1.3300 4.9050 1.3900 ;
      RECT 4.6950 1.2400 4.9050 1.3300 ;
      RECT 4.5150 0.6800 5.5350 0.7700 ;
      RECT 5.4450 0.7700 5.5350 1.2250 ;
      RECT 4.5150 1.4700 4.7250 1.5600 ;
      RECT 4.5150 0.7700 4.6050 1.4700 ;
  END
END MXIT4_X1M_A12TH

MACRO MXIT4_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.3850 0.3200 0.5550 0.3900 ;
        RECT 2.0450 0.3200 2.1350 0.6900 ;
        RECT 3.4800 0.3200 3.6500 0.3800 ;
        RECT 4.0600 0.3200 4.2300 0.3900 ;
        RECT 5.4550 0.3200 5.6250 0.5600 ;
        RECT 6.0300 0.3200 6.1200 0.8850 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1800 0.5500 1.3900 ;
        RECT 0.4500 0.9900 0.5900 1.1800 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3600 1.2200 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.1700 3.5500 1.6050 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 1.0500 2.4350 1.1500 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END D

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 0.8500 2.5550 0.9500 ;
        RECT 1.7950 0.9500 1.8950 1.1600 ;
    END
    ANTENNAGATEAREA 0.1818 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9350 1.0500 5.4500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END S1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.3500 5.8500 1.5050 ;
        RECT 5.6500 1.5050 5.8450 1.5900 ;
        RECT 5.7500 0.6850 5.8500 1.3500 ;
        RECT 5.7550 1.5900 5.8450 1.7400 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 3.4800 2.0300 3.6500 2.0800 ;
        RECT 2.0050 2.0250 2.1750 2.0800 ;
        RECT 4.0450 2.0250 4.2150 2.0800 ;
        RECT 0.3450 1.8650 0.4350 2.0800 ;
        RECT 5.4350 1.5000 5.5250 2.0800 ;
        RECT 6.0300 1.4950 6.1200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5250 1.8150 1.1050 1.9050 ;
      RECT 0.5250 1.7550 0.6150 1.8150 ;
      RECT 0.0600 1.6650 0.6150 1.7550 ;
      RECT 0.0600 0.4800 1.6650 0.5700 ;
      RECT 0.0600 1.3750 0.1750 1.6650 ;
      RECT 0.0600 0.5700 0.1500 1.3750 ;
      RECT 1.2550 1.8150 1.6750 1.9050 ;
      RECT 1.2550 1.7250 1.3450 1.8150 ;
      RECT 0.7050 1.6350 1.3450 1.7250 ;
      RECT 0.7050 0.7550 0.7950 1.6350 ;
      RECT 0.6250 0.6650 1.1000 0.7550 ;
      RECT 2.3200 1.3300 2.4100 1.5350 ;
      RECT 2.3200 1.2400 2.7600 1.3300 ;
      RECT 2.6700 0.7500 2.7600 1.2400 ;
      RECT 2.3200 0.6600 2.7600 0.7500 ;
      RECT 2.3200 0.5400 2.4100 0.6600 ;
      RECT 2.0750 1.6500 2.5900 1.7400 ;
      RECT 2.0750 1.5400 2.1650 1.6500 ;
      RECT 2.5000 1.5200 2.5900 1.6500 ;
      RECT 1.7750 1.4500 2.1650 1.5400 ;
      RECT 2.5000 1.4300 2.9600 1.5200 ;
      RECT 2.8700 0.8500 2.9600 1.4300 ;
      RECT 1.7750 1.3550 1.8650 1.4500 ;
      RECT 1.5800 1.2650 1.8650 1.3550 ;
      RECT 1.5800 0.6600 1.8650 0.7500 ;
      RECT 1.7750 0.4800 1.8650 0.6600 ;
      RECT 1.5800 1.2350 1.6700 1.2650 ;
      RECT 1.1150 1.1450 1.6700 1.2350 ;
      RECT 1.5800 0.7500 1.6700 1.1450 ;
      RECT 3.2300 0.6800 3.3200 1.7000 ;
      RECT 2.5850 0.4800 3.7000 0.5700 ;
      RECT 3.6100 0.5700 3.7000 1.0900 ;
      RECT 2.6800 1.6300 3.1400 1.7200 ;
      RECT 3.0500 0.5700 3.1400 1.6300 ;
      RECT 1.8750 1.8300 4.0600 1.9200 ;
      RECT 3.9700 1.0850 4.0600 1.8300 ;
      RECT 1.8750 1.7250 1.9650 1.8300 ;
      RECT 1.5000 1.6350 1.9650 1.7250 ;
      RECT 1.5000 1.5450 1.5900 1.6350 ;
      RECT 0.9150 1.4550 1.5900 1.5450 ;
      RECT 0.9150 1.0350 1.0050 1.4550 ;
      RECT 0.9150 0.9450 1.3000 1.0350 ;
      RECT 1.2100 0.7550 1.3000 0.9450 ;
      RECT 1.2100 0.6650 1.4100 0.7550 ;
      RECT 4.3600 0.6800 4.4500 1.6150 ;
      RECT 4.1600 1.7800 4.9900 1.8700 ;
      RECT 4.9000 1.4400 4.9900 1.7800 ;
      RECT 3.7900 0.4800 5.0450 0.5700 ;
      RECT 4.1600 0.5700 4.2500 1.7800 ;
      RECT 3.7900 0.5700 3.8800 1.6200 ;
      RECT 5.1650 1.3300 5.2550 1.5000 ;
      RECT 4.7350 1.2400 5.2550 1.3300 ;
      RECT 4.7350 0.8500 5.3150 0.9400 ;
      RECT 4.7350 0.9400 4.8250 1.2400 ;
      RECT 4.5550 0.6700 5.6600 0.7600 ;
      RECT 5.5700 0.7600 5.6600 1.2100 ;
      RECT 4.5550 1.4650 4.7800 1.5550 ;
      RECT 4.5550 0.7600 4.6450 1.4650 ;
  END
END MXIT4_X1P4M_A12TH

MACRO MXIT4_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 1.8950 0.3200 1.9850 0.6650 ;
        RECT 3.0700 0.3200 3.2800 0.3700 ;
        RECT 3.6300 0.3200 3.8400 0.3850 ;
        RECT 4.1700 0.3200 4.3800 0.3850 ;
        RECT 5.4550 0.3200 5.6250 0.4000 ;
        RECT 6.0250 0.3200 6.1250 0.6700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7700 1.4100 5.9500 1.7200 ;
        RECT 5.7700 0.5250 5.8700 1.4100 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9700 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.087 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8000 0.3500 1.2200 ;
    END
    ANTENNAGATEAREA 0.087 ;
  END B

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8850 1.0500 5.2550 1.1750 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END S1

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.7100 3.1500 1.1650 ;
    END
    ANTENNAGATEAREA 0.087 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7450 1.0400 2.1200 1.1550 ;
    END
    ANTENNAGATEAREA 0.087 ;
  END D

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5350 0.8500 2.3700 0.9500 ;
        RECT 1.5350 0.9500 1.6350 1.1550 ;
        RECT 2.2800 0.9500 2.3700 1.1100 ;
    END
    ANTENNAGATEAREA 0.2151 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 4.2300 2.0200 4.3200 2.0800 ;
        RECT 3.6900 2.0100 3.7800 2.0800 ;
        RECT 0.3050 2.0050 0.4900 2.0800 ;
        RECT 6.0250 1.7700 6.1250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0450 1.8150 1.0050 1.9050 ;
      RECT 0.0450 0.5100 1.2650 0.5700 ;
      RECT 0.0450 0.4800 1.5150 0.5100 ;
      RECT 1.1750 0.4200 1.5150 0.4800 ;
      RECT 0.0450 1.4950 0.1750 1.8150 ;
      RECT 0.0450 0.5700 0.1350 1.4950 ;
      RECT 1.1700 1.8700 1.5400 1.9600 ;
      RECT 1.1700 1.7250 1.2600 1.8700 ;
      RECT 0.6500 1.6350 1.2600 1.7250 ;
      RECT 0.6500 0.7700 0.7400 1.6350 ;
      RECT 0.5600 0.6800 0.9850 0.7700 ;
      RECT 2.1550 1.2450 2.5500 1.3350 ;
      RECT 2.4600 0.7550 2.5500 1.2450 ;
      RECT 2.1700 0.6650 2.5500 0.7550 ;
      RECT 2.1550 1.3350 2.2450 1.5350 ;
      RECT 2.1700 0.5150 2.2600 0.6650 ;
      RECT 1.9250 1.6500 2.4250 1.7400 ;
      RECT 2.3350 1.5150 2.4250 1.6500 ;
      RECT 2.3350 1.4250 2.7500 1.5150 ;
      RECT 2.6600 0.9200 2.7500 1.4250 ;
      RECT 1.9250 1.5700 2.0150 1.6500 ;
      RECT 1.6250 1.4800 2.0150 1.5700 ;
      RECT 1.3350 1.2350 1.4250 1.2650 ;
      RECT 1.0100 1.1450 1.4250 1.2350 ;
      RECT 1.3350 0.7500 1.4250 1.1450 ;
      RECT 1.6250 1.3550 1.7150 1.4800 ;
      RECT 1.3350 1.2650 1.7150 1.3550 ;
      RECT 1.3350 0.6600 1.7150 0.7500 ;
      RECT 1.6250 0.5650 1.7150 0.6600 ;
      RECT 2.8400 0.6800 2.9300 1.5150 ;
      RECT 1.7250 1.8300 3.2900 1.9200 ;
      RECT 3.2000 1.7200 3.2900 1.8300 ;
      RECT 3.2000 1.6300 3.5100 1.7200 ;
      RECT 3.4200 1.2050 3.5100 1.6300 ;
      RECT 1.3950 1.5450 1.4850 1.6800 ;
      RECT 0.8300 1.4550 1.4850 1.5450 ;
      RECT 0.8300 1.0350 0.9200 1.4550 ;
      RECT 0.8300 0.9450 1.1650 1.0350 ;
      RECT 1.0750 0.7700 1.1650 0.9450 ;
      RECT 1.0750 0.6800 1.2450 0.7700 ;
      RECT 1.7250 1.7700 1.8150 1.8300 ;
      RECT 1.3950 1.6800 1.8150 1.7700 ;
      RECT 2.5250 1.6250 3.1100 1.7150 ;
      RECT 3.0200 1.4800 3.1100 1.6250 ;
      RECT 3.0200 1.3900 3.3300 1.4800 ;
      RECT 3.2400 0.5700 3.3300 1.3900 ;
      RECT 2.4300 0.4800 3.8700 0.5700 ;
      RECT 3.7800 0.5700 3.8700 1.0400 ;
      RECT 3.7800 1.0400 3.9450 1.2100 ;
      RECT 4.4900 1.6500 5.1400 1.7400 ;
      RECT 3.3800 1.8300 4.5800 1.9200 ;
      RECT 4.4900 1.7400 4.5800 1.8300 ;
      RECT 3.6000 0.8500 3.6900 1.8300 ;
      RECT 3.4200 0.7600 3.6900 0.8500 ;
      RECT 4.7200 1.3700 4.8100 1.6500 ;
      RECT 3.4200 0.6800 3.5100 0.7600 ;
      RECT 4.4800 1.2800 4.8100 1.3700 ;
      RECT 4.4800 0.6600 4.5700 1.2800 ;
      RECT 3.9600 0.4800 5.1600 0.5700 ;
      RECT 3.9600 1.5700 4.1250 1.7400 ;
      RECT 4.0350 1.5500 4.1250 1.5700 ;
      RECT 4.0350 1.4600 4.6100 1.5500 ;
      RECT 4.0350 0.7600 4.1250 1.4600 ;
      RECT 3.9600 0.5700 4.1250 0.7600 ;
      RECT 5.2100 1.4850 5.4450 1.5750 ;
      RECT 5.3550 0.9300 5.4450 1.4850 ;
      RECT 4.6600 0.8400 5.4450 0.9300 ;
      RECT 4.6600 0.9300 4.7500 1.1700 ;
      RECT 4.6900 1.8300 5.6800 1.9200 ;
      RECT 5.5900 0.7500 5.6800 1.8300 ;
      RECT 4.6850 0.6600 5.6800 0.7500 ;
  END
END MXIT4_X2M_A12TH

MACRO MXIT4_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 0.2450 0.3200 0.3450 0.6700 ;
        RECT 4.9250 0.3200 5.0150 0.8450 ;
        RECT 5.4750 0.3200 5.5650 0.5750 ;
        RECT 6.0150 0.3200 6.1050 0.5900 ;
        RECT 8.3000 0.3200 8.5100 0.3600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 0.5750 2.0300 0.7850 2.0800 ;
        RECT 2.7600 2.0250 2.9300 2.0800 ;
        RECT 3.2800 2.0250 3.4500 2.0800 ;
        RECT 1.7000 1.8350 1.7900 2.0800 ;
        RECT 2.2450 1.8350 2.3350 2.0800 ;
        RECT 7.8350 1.8300 7.9350 2.0800 ;
        RECT 8.3550 1.7700 8.4550 2.0800 ;
        RECT 0.0850 1.7100 0.1750 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0900 0.8500 8.7100 0.9500 ;
        RECT 8.6100 0.9500 8.7100 1.3000 ;
        RECT 8.6200 0.5300 8.7100 0.8500 ;
        RECT 8.0900 0.5200 8.1900 0.8500 ;
        RECT 8.0950 1.3000 8.7100 1.4000 ;
        RECT 8.0950 1.4000 8.1950 1.7400 ;
        RECT 8.6200 1.4000 8.7100 1.7400 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7700 1.0500 3.1900 1.1500 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.9400 4.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END D

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.3500 1.0500 7.7700 1.1500 ;
    END
    ANTENNAGATEAREA 0.186 ;
  END S1

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0000 0.3750 1.4700 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5050 0.8500 2.3900 0.9500 ;
        RECT 1.5050 0.9500 1.5950 1.0950 ;
        RECT 2.3000 0.9500 2.3900 1.0500 ;
        RECT 2.3000 0.5700 2.3900 0.8500 ;
        RECT 1.3000 1.0950 1.5950 1.1850 ;
        RECT 2.3000 1.0500 2.4700 1.1500 ;
        RECT 2.3000 0.4800 4.2450 0.5700 ;
        RECT 4.1550 0.5700 4.2450 1.1500 ;
    END
    ANTENNAGATEAREA 0.2682 ;
  END S0

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7050 1.0500 2.1900 1.1500 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.8250 1.4550 2.1250 1.5450 ;
      RECT 1.3250 0.6300 2.0500 0.7200 ;
      RECT 1.8800 0.4300 2.0500 0.6300 ;
      RECT 1.3950 0.4300 1.5650 0.6300 ;
      RECT 0.8250 0.9600 0.9150 1.4550 ;
      RECT 0.8250 0.8700 1.4150 0.9600 ;
      RECT 1.3250 0.7200 1.4150 0.8700 ;
      RECT 3.0000 1.6200 3.6850 1.7100 ;
      RECT 3.5950 1.1350 3.6850 1.6200 ;
      RECT 3.4100 1.0450 3.6850 1.1350 ;
      RECT 3.4100 0.9350 3.5000 1.0450 ;
      RECT 3.2600 0.8450 3.5000 0.9350 ;
      RECT 1.0700 1.2750 3.4850 1.3650 ;
      RECT 3.3950 1.3650 3.4850 1.4850 ;
      RECT 2.5200 0.6650 4.0650 0.7550 ;
      RECT 3.9750 0.7550 4.0650 1.2600 ;
      RECT 3.9750 1.2600 4.1500 1.3500 ;
      RECT 2.4800 1.3650 2.6600 1.5250 ;
      RECT 2.5700 0.9300 2.6600 1.2750 ;
      RECT 2.5200 0.7550 2.6600 0.9300 ;
      RECT 1.0700 1.0650 1.1600 1.2750 ;
      RECT 4.0600 1.4700 4.8100 1.5600 ;
      RECT 4.3350 0.7250 4.6750 0.8150 ;
      RECT 4.5850 0.4150 4.6750 0.7250 ;
      RECT 4.3350 0.8150 4.4250 1.4700 ;
      RECT 4.3350 0.4850 4.4250 0.7250 ;
      RECT 3.7750 1.6500 5.1050 1.7400 ;
      RECT 5.0150 1.0250 5.1050 1.6500 ;
      RECT 3.7750 0.9350 3.8650 1.6500 ;
      RECT 3.6750 0.8450 3.8650 0.9350 ;
      RECT 2.7850 1.8300 5.6300 1.9200 ;
      RECT 5.5400 1.0300 5.6300 1.8300 ;
      RECT 2.7850 1.7250 2.8750 1.8300 ;
      RECT 0.6450 1.6350 2.8750 1.7250 ;
      RECT 0.6450 0.7800 0.7350 1.6350 ;
      RECT 0.6450 0.6900 1.2350 0.7800 ;
      RECT 1.1450 0.4100 1.2350 0.6900 ;
      RECT 5.7400 1.8300 7.1750 1.9200 ;
      RECT 5.7400 0.9550 5.8300 1.8300 ;
      RECT 5.6800 0.8650 6.6750 0.9550 ;
      RECT 6.2200 1.4500 6.6750 1.5400 ;
      RECT 6.2200 1.1400 6.3100 1.4500 ;
      RECT 6.2200 1.0500 6.8850 1.1400 ;
      RECT 6.7950 0.7750 6.8850 1.0500 ;
      RECT 5.2000 0.6850 7.1950 0.7750 ;
      RECT 5.2000 0.7750 5.2900 1.7100 ;
      RECT 5.2000 0.5650 5.2900 0.6850 ;
      RECT 7.5550 1.3950 7.6450 1.5150 ;
      RECT 7.1500 1.3400 7.6450 1.3950 ;
      RECT 6.4200 1.3050 7.6450 1.3400 ;
      RECT 7.1500 0.8700 7.6450 0.9600 ;
      RECT 7.5550 0.7500 7.6450 0.8700 ;
      RECT 6.4200 1.2500 7.2400 1.3050 ;
      RECT 7.1500 0.9600 7.2400 1.2500 ;
      RECT 7.8800 1.0850 8.4000 1.1750 ;
      RECT 7.2650 1.7200 7.4350 1.9600 ;
      RECT 6.2050 1.6300 7.9700 1.7200 ;
      RECT 7.8800 1.1750 7.9700 1.6300 ;
      RECT 7.8800 0.5950 7.9700 1.0850 ;
      RECT 6.2150 0.5050 7.9700 0.5950 ;
      RECT 0.3600 1.8300 1.5650 1.9200 ;
      RECT 0.3600 1.9200 0.4500 1.9900 ;
      RECT 0.3600 1.6700 0.4500 1.8300 ;
      RECT 0.3600 1.5800 0.5550 1.6700 ;
      RECT 0.4650 0.5750 0.5550 1.5800 ;
      RECT 0.4650 0.4850 1.0350 0.5750 ;
  END
END MXIT4_X3M_A12TH

MACRO MXT2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.4200 0.3200 0.5900 0.3600 ;
        RECT 1.7500 0.3200 1.8500 0.7350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6050 0.9150 1.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0333 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0300 0.5700 1.4150 ;
    END
    ANTENNAGATEAREA 0.0333 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9250 0.3500 1.3700 ;
        RECT 0.2500 0.8350 0.5500 0.9250 ;
        RECT 0.4500 0.5700 0.5500 0.8350 ;
        RECT 0.4500 0.4800 1.3350 0.5700 ;
        RECT 1.2450 0.5700 1.3350 1.4700 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0300 1.5700 2.1500 1.9850 ;
        RECT 2.0500 0.9000 2.1500 1.5700 ;
        RECT 2.0150 0.5000 2.1500 0.9000 ;
    END
    ANTENNADIFFAREA 0.14175 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6950 0.6700 0.7850 1.7200 ;
      RECT 0.0500 1.8300 0.9650 1.9200 ;
      RECT 0.8750 1.1750 0.9650 1.8300 ;
      RECT 0.0500 1.6600 0.1850 1.8300 ;
      RECT 0.0500 0.7900 0.1400 1.6600 ;
      RECT 0.0500 0.6050 0.1700 0.7900 ;
      RECT 1.3000 1.5800 1.5150 1.6700 ;
      RECT 1.4250 0.6600 1.5150 1.5800 ;
      RECT 1.0550 1.7850 1.9400 1.8750 ;
      RECT 1.8500 1.0600 1.9400 1.7850 ;
      RECT 1.0550 0.8300 1.1450 1.7850 ;
      RECT 0.8950 0.7400 1.1450 0.8300 ;
  END
END MXT2_X0P5M_A12TH

MACRO MXT2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.4100 0.3200 0.5800 0.3900 ;
        RECT 1.7700 0.3200 1.8700 0.8100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6200 0.9500 1.7500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5700 1.4300 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9200 0.3500 1.4550 ;
        RECT 0.2500 0.8300 0.5450 0.9200 ;
        RECT 0.4550 0.5700 0.5450 0.8300 ;
        RECT 0.4550 0.4800 1.3450 0.5700 ;
        RECT 1.2550 0.5700 1.3450 1.5350 ;
        RECT 0.7900 0.4450 0.9600 0.4800 ;
    END
    ANTENNAGATEAREA 0.0774 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0300 1.5250 2.1500 1.9300 ;
        RECT 2.0500 0.9200 2.1500 1.5250 ;
        RECT 2.0150 0.5100 2.1500 0.9200 ;
    END
    ANTENNADIFFAREA 0.1816 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.6950 2.0350 1.9050 2.0800 ;
        RECT 0.3600 1.9600 0.4600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6150 1.5500 0.7850 1.6400 ;
      RECT 0.6950 0.7300 0.7850 1.5500 ;
      RECT 0.0500 1.7500 0.9750 1.8400 ;
      RECT 0.8850 1.2050 0.9750 1.7500 ;
      RECT 0.0500 1.6500 0.1700 1.7500 ;
      RECT 0.0500 0.7800 0.1400 1.6500 ;
      RECT 0.0500 0.5900 0.1700 0.7800 ;
      RECT 1.3200 1.6450 1.5250 1.7350 ;
      RECT 1.4350 0.7100 1.5250 1.6450 ;
      RECT 1.0650 1.8300 1.9400 1.9200 ;
      RECT 1.8500 1.0450 1.9400 1.8300 ;
      RECT 1.0650 0.8700 1.1550 1.8300 ;
      RECT 0.8950 0.7800 1.1550 0.8700 ;
  END
END MXT2_X0P7M_A12TH

MACRO MXT2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.3700 ;
        RECT 1.7700 0.3200 1.8600 0.6250 ;
    END
  END VSS

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8900 0.3600 1.2650 ;
        RECT 0.2500 0.8000 0.5450 0.8900 ;
        RECT 0.4550 0.5700 0.5450 0.8000 ;
        RECT 0.4550 0.4800 1.3700 0.5700 ;
        RECT 0.9050 0.5700 0.9950 1.0650 ;
        RECT 1.2800 0.5700 1.3700 1.4850 ;
    END
    ANTENNAGATEAREA 0.1002 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6400 1.2100 1.7500 1.6300 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1650 0.5500 1.3900 ;
        RECT 0.4500 0.9900 0.5900 1.1650 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0300 1.2900 2.1500 1.7450 ;
        RECT 2.0500 0.9150 2.1500 1.2900 ;
        RECT 2.0300 0.5300 2.1500 0.9150 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7050 0.6600 0.7950 1.7150 ;
      RECT 0.0600 1.8250 0.9950 1.9150 ;
      RECT 0.9050 1.1750 0.9950 1.8250 ;
      RECT 0.0600 1.4900 0.1750 1.8250 ;
      RECT 0.0600 0.7300 0.1500 1.4900 ;
      RECT 0.0600 0.5150 0.1750 0.7300 ;
      RECT 1.3000 1.6100 1.5500 1.7000 ;
      RECT 1.4600 0.4400 1.5500 1.6100 ;
      RECT 1.1000 1.8300 1.9350 1.9200 ;
      RECT 1.8450 1.0400 1.9350 1.8300 ;
      RECT 1.1000 0.6800 1.1900 1.8300 ;
  END
END MXT2_X1M_A12TH

MACRO MXT2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.2950 0.3200 0.4850 0.3900 ;
        RECT 1.6950 0.3200 1.7950 0.7150 ;
        RECT 2.2250 0.3200 2.3250 0.7250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2150 0.5500 1.3900 ;
        RECT 0.4500 0.9900 0.5900 1.2150 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9000 0.3600 1.3350 ;
        RECT 0.2500 0.8000 0.5500 0.9000 ;
        RECT 0.4500 0.5800 0.5500 0.8000 ;
        RECT 0.4500 0.4800 1.3500 0.5800 ;
        RECT 0.8800 0.5800 0.9700 1.0650 ;
        RECT 1.2500 0.5800 1.3500 1.4800 ;
    END
    ANTENNAGATEAREA 0.1323 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6300 0.8100 1.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9000 2.1500 1.5000 ;
        RECT 1.9700 1.5000 2.1500 1.6000 ;
        RECT 1.9700 0.8000 2.1500 0.9000 ;
        RECT 1.9700 1.6000 2.0700 1.9250 ;
        RECT 1.9700 0.4200 2.0700 0.8000 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.6500 2.0450 1.8400 2.0800 ;
        RECT 2.2250 1.6850 2.3250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6900 0.6900 0.7800 1.7000 ;
      RECT 0.0450 1.8250 0.9700 1.9150 ;
      RECT 0.8800 1.1750 0.9700 1.8250 ;
      RECT 0.0450 1.5000 0.1750 1.8250 ;
      RECT 0.0450 0.7000 0.1350 1.5000 ;
      RECT 0.0450 0.6100 0.2350 0.7000 ;
      RECT 1.4400 0.4300 1.5300 1.7200 ;
      RECT 1.0600 1.8300 1.7450 1.9200 ;
      RECT 1.6550 1.3900 1.7450 1.8300 ;
      RECT 1.6550 1.3000 1.9400 1.3900 ;
      RECT 1.0600 0.6900 1.1500 1.8300 ;
  END
END MXT2_X1P4M_A12TH

MACRO MXT2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 1.6950 0.3200 1.7950 0.6400 ;
        RECT 2.2250 0.3200 2.3250 0.6400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9000 2.3500 1.5350 ;
        RECT 1.9700 1.5350 2.3500 1.6350 ;
        RECT 1.9700 0.8000 2.3500 0.9000 ;
        RECT 1.9700 1.6350 2.0700 1.9550 ;
        RECT 1.9700 0.4750 2.0700 0.8000 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6300 0.8100 1.7500 1.2150 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1650 0.5500 1.3900 ;
        RECT 0.4500 0.9900 0.5900 1.1650 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8900 0.3600 1.2800 ;
        RECT 0.2500 0.7900 0.5500 0.8900 ;
        RECT 0.4500 0.5700 0.5500 0.7900 ;
        RECT 0.4500 0.4800 1.3500 0.5700 ;
        RECT 0.8900 0.5700 0.9800 1.0700 ;
        RECT 1.2500 0.5700 1.3500 1.4800 ;
    END
    ANTENNAGATEAREA 0.177 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 2.2250 1.7700 2.3250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6850 0.6850 0.7750 1.7150 ;
      RECT 0.0600 1.8250 0.9800 1.9150 ;
      RECT 0.8900 1.1800 0.9800 1.8250 ;
      RECT 0.0600 1.4700 0.1750 1.8250 ;
      RECT 0.0600 0.7050 0.1500 1.4700 ;
      RECT 0.0600 0.4950 0.1750 0.7050 ;
      RECT 1.2800 1.6100 1.5300 1.7000 ;
      RECT 1.4400 0.4400 1.5300 1.6100 ;
      RECT 1.6400 1.3250 2.1350 1.4150 ;
      RECT 2.0450 1.0200 2.1350 1.3250 ;
      RECT 1.0700 1.8300 1.7300 1.9200 ;
      RECT 1.6400 1.4150 1.7300 1.8300 ;
      RECT 1.0700 0.6850 1.1600 1.8300 ;
  END
END MXT2_X2M_A12TH

MACRO MXT2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.8300 ;
        RECT 0.5900 0.3200 0.7400 0.5650 ;
        RECT 1.1200 0.3200 1.2500 0.5750 ;
        RECT 2.6700 0.3200 2.8400 0.5550 ;
        RECT 3.2100 0.3200 3.3800 0.5700 ;
        RECT 3.7650 0.3200 3.8650 0.6800 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3750 1.3900 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9850 1.0500 1.6550 1.1500 ;
    END
    ANTENNAGATEAREA 0.2592 ;
  END S0

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7600 1.0500 3.2000 1.1700 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.9500 4.1500 1.2500 ;
        RECT 3.5050 1.2500 4.1500 1.3500 ;
        RECT 3.5050 0.8500 4.1500 0.9500 ;
        RECT 3.5050 1.3500 3.6050 1.7300 ;
        RECT 4.0250 1.3500 4.1250 1.7250 ;
        RECT 4.0250 0.5150 4.1250 0.8500 ;
        RECT 3.5050 0.5100 3.6050 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 3.2100 1.8400 3.3800 2.0800 ;
        RECT 1.1350 1.8350 1.2350 2.0800 ;
        RECT 0.6150 1.8000 0.7150 2.0800 ;
        RECT 2.7200 1.7550 2.8100 2.0800 ;
        RECT 3.7650 1.7550 3.8650 2.0800 ;
        RECT 0.0950 1.5650 0.1950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 1.6100 1.8100 1.7000 ;
      RECT 0.3550 0.6650 2.3500 0.7550 ;
      RECT 0.3550 1.7000 0.4550 1.9800 ;
      RECT 0.3550 0.4200 0.4550 0.6650 ;
      RECT 0.5800 0.7900 0.6700 1.6100 ;
      RECT 0.3550 0.7550 0.6700 0.7900 ;
      RECT 0.7600 1.4000 1.9900 1.4900 ;
      RECT 1.9000 1.1500 1.9900 1.4000 ;
      RECT 1.9000 1.0500 2.3750 1.1500 ;
      RECT 0.7600 0.8450 1.0300 0.9350 ;
      RECT 0.7600 0.9350 0.8500 1.4000 ;
      RECT 2.2000 1.3250 3.1300 1.4150 ;
      RECT 1.6100 0.8450 3.1300 0.9350 ;
      RECT 2.2000 1.4150 2.2900 1.6800 ;
      RECT 2.4650 0.9350 2.5550 1.3250 ;
      RECT 3.3000 1.0500 3.8300 1.1500 ;
      RECT 1.3450 1.7900 2.6100 1.8800 ;
      RECT 2.5200 1.6200 2.6100 1.7900 ;
      RECT 2.4600 0.5700 2.5500 0.6650 ;
      RECT 1.3600 0.4800 2.5500 0.5700 ;
      RECT 2.5200 1.5300 3.3900 1.6200 ;
      RECT 3.3000 1.1500 3.3900 1.5300 ;
      RECT 3.3000 0.7550 3.3900 1.0500 ;
      RECT 2.4600 0.6650 3.3900 0.7550 ;
  END
END MXT2_X3M_A12TH

MACRO MXT2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6900 ;
        RECT 0.5600 0.3200 0.7300 0.5450 ;
        RECT 1.1150 0.3200 1.2150 0.4500 ;
        RECT 2.6550 0.3200 2.7550 0.5500 ;
        RECT 3.1500 0.3200 3.3200 0.5700 ;
        RECT 3.7050 0.3200 3.8050 0.6900 ;
        RECT 4.2250 0.3200 4.3250 0.6900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0100 0.3550 1.3900 ;
    END
    ANTENNAGATEAREA 0.1734 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9600 1.0500 1.6300 1.1500 ;
    END
    ANTENNAGATEAREA 0.3372 ;
  END S0

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6950 1.0500 3.1450 1.1700 ;
    END
    ANTENNAGATEAREA 0.1734 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.9500 4.1500 1.2500 ;
        RECT 3.4450 1.2500 4.1500 1.3500 ;
        RECT 3.4450 0.8500 4.1500 0.9500 ;
        RECT 3.4450 1.3500 3.5450 1.7300 ;
        RECT 3.9650 1.3500 4.0650 1.7250 ;
        RECT 3.9650 0.5150 4.0650 0.8500 ;
        RECT 3.4450 0.5000 3.5450 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 2.6600 1.9000 2.7500 2.0800 ;
        RECT 3.1500 1.8400 3.3200 2.0800 ;
        RECT 1.1150 1.8200 1.2150 2.0800 ;
        RECT 0.5950 1.8000 0.6950 2.0800 ;
        RECT 3.7050 1.7550 3.8050 2.0800 ;
        RECT 4.2250 1.7550 4.3250 2.0800 ;
        RECT 0.0750 1.6900 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7400 1.4000 1.9450 1.4900 ;
      RECT 1.8550 1.1500 1.9450 1.4000 ;
      RECT 1.8550 1.0500 2.3000 1.1500 ;
      RECT 0.7400 0.8450 1.0300 0.9350 ;
      RECT 0.7400 0.9350 0.8300 1.4000 ;
      RECT 0.3350 1.6100 1.7800 1.7000 ;
      RECT 0.3000 0.6650 2.3000 0.7550 ;
      RECT 0.5600 0.7550 0.6500 1.6100 ;
      RECT 0.3350 1.7000 0.4350 1.9800 ;
      RECT 0.3000 0.4650 0.4700 0.6650 ;
      RECT 2.1100 1.4400 3.0700 1.5300 ;
      RECT 1.5700 0.8450 3.0700 0.9350 ;
      RECT 2.1100 1.5300 2.2800 1.7050 ;
      RECT 2.1100 1.4150 2.5000 1.4400 ;
      RECT 2.4100 0.9350 2.5000 1.4150 ;
      RECT 3.2450 1.0500 3.7700 1.1500 ;
      RECT 1.3250 1.8300 2.5000 1.9200 ;
      RECT 2.4100 1.7350 2.5000 1.8300 ;
      RECT 2.4100 0.5700 2.5000 0.6650 ;
      RECT 1.3250 0.4800 2.5000 0.5700 ;
      RECT 2.4100 1.6450 3.3350 1.7350 ;
      RECT 3.2450 1.1500 3.3350 1.6450 ;
      RECT 3.2450 0.7550 3.3350 1.0500 ;
      RECT 2.4100 0.6650 3.3350 0.7550 ;
  END
END MXT2_X4M_A12TH

MACRO MXT2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6750 ;
        RECT 0.8100 0.3200 1.0000 0.5700 ;
        RECT 1.3450 0.3200 1.5350 0.5700 ;
        RECT 3.9850 0.3200 4.1350 0.5650 ;
        RECT 4.5350 0.3200 4.6950 0.5650 ;
        RECT 5.1050 0.3200 5.2050 0.6800 ;
        RECT 5.6450 0.3200 5.7450 0.6800 ;
        RECT 6.1850 0.3200 6.2850 0.6800 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2950 1.0500 0.7350 1.1500 ;
    END
    ANTENNAGATEAREA 0.2529 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 1.0500 2.3250 1.1500 ;
    END
    ANTENNAGATEAREA 0.4959 ;
  END S0

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9650 1.0500 4.4500 1.1700 ;
    END
    ANTENNAGATEAREA 0.2529 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.9500 6.1500 1.2500 ;
        RECT 4.8450 1.2500 6.1500 1.3500 ;
        RECT 4.8450 0.8500 6.1500 0.9500 ;
        RECT 4.8450 1.3500 4.9450 1.7300 ;
        RECT 5.3850 1.3500 5.4850 1.7250 ;
        RECT 5.9250 1.3500 6.0250 1.7250 ;
        RECT 5.3850 0.5150 5.4850 0.8500 ;
        RECT 5.9250 0.5150 6.0250 0.8500 ;
        RECT 4.8450 0.5100 4.9450 0.8500 ;
    END
    ANTENNADIFFAREA 1.0075 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.8200 1.9300 0.9900 2.0800 ;
        RECT 1.3450 1.8650 1.5350 2.0800 ;
        RECT 3.9650 1.8050 4.1550 2.0800 ;
        RECT 4.5150 1.8050 4.7100 2.0800 ;
        RECT 5.1050 1.7550 5.2050 2.0800 ;
        RECT 5.6450 1.7550 5.7450 2.0800 ;
        RECT 6.1850 1.7550 6.2850 2.0800 ;
        RECT 0.3350 1.7000 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0750 1.4500 2.9400 1.5400 ;
      RECT 2.8500 1.1500 2.9400 1.4500 ;
      RECT 2.8500 1.0500 3.3000 1.1500 ;
      RECT 1.0750 0.8450 1.7950 0.9350 ;
      RECT 1.0750 0.9350 1.1650 1.4500 ;
      RECT 0.8800 1.6500 2.6150 1.7400 ;
      RECT 0.8800 0.6650 3.6550 0.7550 ;
      RECT 0.0750 1.5900 0.1750 1.9450 ;
      RECT 0.0800 0.4200 0.1800 0.8000 ;
      RECT 0.5950 1.5900 0.6950 1.9450 ;
      RECT 0.5950 0.4200 0.6950 0.8000 ;
      RECT 0.8800 1.5900 0.9700 1.6500 ;
      RECT 0.0750 1.5000 0.9700 1.5900 ;
      RECT 0.8800 0.8900 0.9700 1.5000 ;
      RECT 0.0800 0.8000 0.9700 0.8900 ;
      RECT 0.8800 0.7550 0.9700 0.8000 ;
      RECT 3.5050 1.3250 4.4450 1.4150 ;
      RECT 1.9050 0.8450 4.4450 0.9350 ;
      RECT 2.9200 1.6500 3.5950 1.7400 ;
      RECT 3.5050 1.4150 3.5950 1.6500 ;
      RECT 3.5050 0.9350 3.5950 1.3250 ;
      RECT 4.5800 1.0550 5.7650 1.1550 ;
      RECT 2.1450 1.8300 3.8250 1.9200 ;
      RECT 3.7350 1.6200 3.8250 1.8300 ;
      RECT 3.7650 0.5700 3.8550 0.6650 ;
      RECT 2.1450 0.4800 3.8550 0.5700 ;
      RECT 3.7350 1.5300 4.6700 1.6200 ;
      RECT 4.5800 1.1550 4.6700 1.5300 ;
      RECT 4.5800 0.7550 4.6700 1.0550 ;
      RECT 3.7650 0.6650 4.6700 0.7550 ;
  END
END MXT2_X6M_A12TH

MACRO MXT4_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 1.7450 0.3200 1.8450 0.6700 ;
        RECT 3.2250 0.3200 3.3950 0.3600 ;
        RECT 4.4700 0.3200 4.6400 0.5500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0950 0.5500 1.5150 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0000 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9750 3.1500 1.4000 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8050 1.0500 2.1900 1.1500 ;
        RECT 1.8050 1.1500 1.9400 1.2400 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END D

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 0.8500 2.2200 0.9500 ;
        RECT 1.6000 0.9500 1.6900 1.0600 ;
    END
    ANTENNAGATEAREA 0.117 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0600 4.1500 1.4800 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END S1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.0000 4.9500 1.5200 ;
        RECT 4.8300 1.5200 4.9500 1.9400 ;
        RECT 4.8300 0.5700 4.9500 1.0000 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 3.2300 1.8500 3.3300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5550 1.6250 0.7500 1.7150 ;
      RECT 0.6600 1.3650 0.7500 1.6250 ;
      RECT 0.6600 1.2750 0.8100 1.3650 ;
      RECT 0.7200 0.6600 0.8100 1.2750 ;
      RECT 0.0550 1.8050 1.3100 1.8950 ;
      RECT 0.0550 0.4800 1.3300 0.5700 ;
      RECT 1.2400 0.5700 1.3300 0.7700 ;
      RECT 0.0550 1.5050 0.1700 1.8050 ;
      RECT 0.0550 0.7200 0.1450 1.5050 ;
      RECT 0.0550 0.5700 0.1700 0.7200 ;
      RECT 2.0400 1.3800 2.1300 1.5350 ;
      RECT 2.0400 1.2900 2.4200 1.3800 ;
      RECT 2.3300 0.7500 2.4200 1.2900 ;
      RECT 2.0350 0.6600 2.4200 0.7500 ;
      RECT 2.0350 0.5100 2.1250 0.6600 ;
      RECT 1.6550 1.6450 2.3100 1.7350 ;
      RECT 2.2200 1.5600 2.3100 1.6450 ;
      RECT 2.2200 1.4700 2.6000 1.5600 ;
      RECT 2.5100 0.8100 2.6000 1.4700 ;
      RECT 1.6550 1.5350 1.7450 1.6450 ;
      RECT 1.4200 1.4450 1.7450 1.5350 ;
      RECT 1.4200 0.6250 1.6400 0.7150 ;
      RECT 1.4200 1.2000 1.5100 1.4450 ;
      RECT 1.1600 1.1100 1.5100 1.2000 ;
      RECT 1.4200 0.7150 1.5100 1.1100 ;
      RECT 2.8700 0.6800 2.9600 1.7200 ;
      RECT 3.0500 1.6400 4.1600 1.7300 ;
      RECT 3.9900 1.5950 4.1600 1.6400 ;
      RECT 3.7350 1.3500 3.8250 1.6400 ;
      RECT 3.4200 1.2600 3.8250 1.3500 ;
      RECT 3.4200 0.7500 3.5100 1.2600 ;
      RECT 3.4200 0.6600 3.6150 0.7500 ;
      RECT 1.4550 1.8300 3.1400 1.9200 ;
      RECT 3.0500 1.7300 3.1400 1.8300 ;
      RECT 1.4550 1.7150 1.5450 1.8300 ;
      RECT 0.8600 1.6250 1.5450 1.7150 ;
      RECT 0.9800 0.6600 1.0700 1.6250 ;
      RECT 2.3400 0.4800 4.1900 0.5700 ;
      RECT 3.2400 0.5700 3.3300 1.4600 ;
      RECT 3.2400 1.4600 3.6150 1.5500 ;
      RECT 2.4200 1.6500 2.7800 1.7400 ;
      RECT 2.6900 0.5700 2.7800 1.6500 ;
      RECT 4.2750 1.5100 4.4250 1.7300 ;
      RECT 4.3350 0.9500 4.4250 1.5100 ;
      RECT 3.6000 0.8600 4.4250 0.9500 ;
      RECT 3.6000 0.9500 3.6900 1.1350 ;
      RECT 3.6950 1.8200 4.7050 1.9100 ;
      RECT 4.6150 0.7500 4.7050 1.8200 ;
      RECT 3.7250 0.6600 4.7050 0.7500 ;
  END
END MXT4_X0P5M_A12TH

MACRO MXT4_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 1.6950 0.3200 1.8650 0.5700 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0700 0.5500 1.5250 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9150 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9950 3.1500 1.4400 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8100 1.0500 2.1900 1.1500 ;
        RECT 1.8100 1.1500 1.9400 1.2400 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END D

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5700 0.8500 2.2200 0.9500 ;
    END
    ANTENNAGATEAREA 0.1566 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0600 4.1500 1.4800 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END S1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.0000 4.9500 1.5200 ;
        RECT 4.8250 1.5200 4.9500 1.9400 ;
        RECT 4.8300 0.5700 4.9500 1.0000 ;
    END
    ANTENNADIFFAREA 0.1816 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.2900 2.0000 0.5000 2.0800 ;
        RECT 4.4950 1.9450 4.7050 2.0800 ;
        RECT 3.2350 1.8500 3.3350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5600 1.6150 0.7900 1.7050 ;
      RECT 0.7000 0.8850 0.7900 1.6150 ;
      RECT 0.6650 0.6750 0.7900 0.8850 ;
      RECT 0.0550 1.7950 1.2900 1.8850 ;
      RECT 0.0550 0.4800 1.3550 0.5700 ;
      RECT 0.0550 1.5100 0.1700 1.7950 ;
      RECT 0.0550 0.6650 0.1450 1.5100 ;
      RECT 0.0550 0.5700 0.1700 0.6650 ;
      RECT 2.0400 1.3800 2.1300 1.5200 ;
      RECT 2.0400 1.2900 2.4200 1.3800 ;
      RECT 2.3300 0.7500 2.4200 1.2900 ;
      RECT 2.0350 0.6600 2.4200 0.7500 ;
      RECT 2.0350 0.5100 2.1250 0.6600 ;
      RECT 1.6550 1.6450 2.3100 1.7350 ;
      RECT 2.2200 1.5600 2.3100 1.6450 ;
      RECT 2.2200 1.4700 2.6000 1.5600 ;
      RECT 2.5100 0.8100 2.6000 1.4700 ;
      RECT 1.6550 1.5050 1.7450 1.6450 ;
      RECT 1.3200 1.4150 1.7450 1.5050 ;
      RECT 1.3200 0.6600 1.6500 0.7500 ;
      RECT 1.3200 1.1950 1.4100 1.4150 ;
      RECT 1.1250 1.1050 1.4100 1.1950 ;
      RECT 1.3200 0.7500 1.4100 1.1050 ;
      RECT 2.8700 0.6800 2.9600 1.7200 ;
      RECT 2.3000 0.4800 4.1600 0.5700 ;
      RECT 3.2400 0.5700 3.3300 1.4550 ;
      RECT 3.2400 1.4550 3.6400 1.5450 ;
      RECT 2.4200 1.6500 2.7800 1.7400 ;
      RECT 2.6900 0.5700 2.7800 1.6500 ;
      RECT 3.0500 1.6500 4.1800 1.7400 ;
      RECT 3.7500 1.3450 3.8400 1.6500 ;
      RECT 3.4200 1.2550 3.8400 1.3450 ;
      RECT 3.4200 0.7600 3.5100 1.2550 ;
      RECT 3.4200 0.6700 3.5950 0.7600 ;
      RECT 1.4550 1.8300 3.1400 1.9200 ;
      RECT 3.0500 1.7400 3.1400 1.8300 ;
      RECT 1.4550 1.7050 1.5450 1.8300 ;
      RECT 0.8800 1.6150 1.5450 1.7050 ;
      RECT 0.8800 1.4750 1.0300 1.6150 ;
      RECT 0.9400 0.6750 1.0300 1.4750 ;
      RECT 4.2400 1.4600 4.4300 1.5500 ;
      RECT 4.3400 0.9400 4.4300 1.4600 ;
      RECT 3.6000 0.8500 4.4300 0.9400 ;
      RECT 3.6000 0.9400 3.6900 1.1350 ;
      RECT 3.7000 1.8300 4.3800 1.9200 ;
      RECT 4.2900 1.7500 4.3800 1.8300 ;
      RECT 4.2900 1.6600 4.7050 1.7500 ;
      RECT 4.6150 0.7600 4.7050 1.6600 ;
      RECT 3.7050 0.6700 4.7050 0.7600 ;
  END
END MXT4_X0P7M_A12TH

MACRO MXT4_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 4.7300 0.3200 4.9000 0.5700 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9800 0.5850 1.1950 ;
        RECT 0.4500 1.1950 0.5500 1.4150 ;
    END
    ANTENNAGATEAREA 0.0921 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9700 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0921 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9700 3.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0921 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6100 1.2500 2.0900 1.3500 ;
        RECT 1.9900 1.0600 2.0900 1.2500 ;
    END
    ANTENNAGATEAREA 0.0921 ;
  END D

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 0.8500 2.3800 0.9500 ;
        RECT 1.6000 0.9500 1.7000 1.1150 ;
        RECT 2.2800 0.9500 2.3800 1.0950 ;
    END
    ANTENNAGATEAREA 0.2178 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.0600 4.1650 1.4800 ;
    END
    ANTENNAGATEAREA 0.1122 ;
  END S1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0300 0.5000 5.1500 1.7500 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0700 1.8300 1.5200 1.9200 ;
      RECT 1.0700 1.7200 1.1600 1.8300 ;
      RECT 0.5400 1.6300 1.1600 1.7200 ;
      RECT 0.6750 0.7500 0.7650 1.6300 ;
      RECT 0.5400 0.6600 1.0000 0.7500 ;
      RECT 0.0550 1.8300 0.9800 1.9200 ;
      RECT 0.0550 0.4800 1.5200 0.5700 ;
      RECT 0.0550 1.5000 0.1700 1.8300 ;
      RECT 0.0550 0.6950 0.1450 1.5000 ;
      RECT 0.0550 0.5700 0.1950 0.6950 ;
      RECT 2.2200 1.3250 2.3100 1.5000 ;
      RECT 2.2200 1.2350 2.5600 1.3250 ;
      RECT 2.4700 0.7500 2.5600 1.2350 ;
      RECT 2.1550 0.6600 2.5600 0.7500 ;
      RECT 2.1550 0.4600 2.3250 0.6600 ;
      RECT 1.9750 1.6450 2.4900 1.7350 ;
      RECT 2.4000 1.5050 2.4900 1.6450 ;
      RECT 2.4000 1.4150 2.7500 1.5050 ;
      RECT 2.6600 0.8600 2.7500 1.4150 ;
      RECT 1.4300 1.2950 1.5200 1.4700 ;
      RECT 1.0350 1.2050 1.5200 1.2950 ;
      RECT 1.0350 1.0800 1.1250 1.2050 ;
      RECT 1.3100 0.7500 1.4000 1.2050 ;
      RECT 1.9750 1.5600 2.0650 1.6450 ;
      RECT 1.4300 1.4700 2.0650 1.5600 ;
      RECT 1.3100 0.6600 1.7700 0.7500 ;
      RECT 3.0200 1.5900 3.1100 1.7150 ;
      RECT 3.0200 1.5000 3.3300 1.5900 ;
      RECT 3.2400 0.8500 3.3300 1.5000 ;
      RECT 3.0200 0.7600 3.3300 0.8500 ;
      RECT 3.0200 0.6800 3.1100 0.7600 ;
      RECT 3.4200 1.6500 4.3250 1.7400 ;
      RECT 1.6700 1.8300 3.5100 1.9200 ;
      RECT 3.4200 1.7400 3.5100 1.8300 ;
      RECT 3.8500 1.2650 3.9400 1.6500 ;
      RECT 3.6000 1.1750 3.9400 1.2650 ;
      RECT 3.6000 0.7700 3.6900 1.1750 ;
      RECT 3.6000 0.6800 3.7700 0.7700 ;
      RECT 1.2500 1.5200 1.3400 1.6500 ;
      RECT 0.8550 1.4300 1.3400 1.5200 ;
      RECT 0.8550 0.9450 0.9450 1.4300 ;
      RECT 0.8550 0.8550 1.2000 0.9450 ;
      RECT 1.1100 0.6600 1.2000 0.8550 ;
      RECT 1.6700 1.7400 1.7600 1.8300 ;
      RECT 1.2500 1.6500 1.7600 1.7400 ;
      RECT 2.4850 0.4800 4.3300 0.5700 ;
      RECT 3.4200 0.5700 3.5100 1.3750 ;
      RECT 3.4200 1.3750 3.7400 1.4650 ;
      RECT 3.6500 1.4650 3.7400 1.5600 ;
      RECT 2.5800 1.6300 2.9300 1.7200 ;
      RECT 2.8400 0.5700 2.9300 1.6300 ;
      RECT 4.4350 1.2800 4.5650 1.6500 ;
      RECT 4.4750 0.9500 4.5650 1.2800 ;
      RECT 3.8050 0.8600 4.5650 0.9500 ;
      RECT 3.8050 0.9500 3.8950 1.0850 ;
      RECT 3.8500 1.8300 4.8600 1.9200 ;
      RECT 4.7600 0.7700 4.8600 1.8300 ;
      RECT 3.8800 0.6800 4.8600 0.7700 ;
  END
END MXT4_X1M_A12TH

MACRO MXT4_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.5600 0.3200 0.7300 0.5250 ;
        RECT 2.3950 0.3200 2.4950 0.7050 ;
        RECT 6.4250 0.3200 6.5250 0.7750 ;
    END
  END VSS

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2600 1.0500 5.5900 1.1500 ;
        RECT 5.4900 1.1500 5.5900 1.3500 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END S1

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 1.2500 0.5100 1.3500 ;
    END
    ANTENNAGATEAREA 0.111 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 0.9500 1.5550 ;
    END
    ANTENNAGATEAREA 0.111 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2500 0.9500 6.3500 1.2900 ;
        RECT 6.1700 1.2900 6.3500 1.3900 ;
        RECT 6.1650 0.8500 6.3500 0.9500 ;
        RECT 6.1700 1.3900 6.2700 1.7650 ;
        RECT 6.1650 0.4700 6.2650 0.8500 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.5450 2.0400 0.7350 2.0800 ;
        RECT 1.0700 2.0400 1.2600 2.0800 ;
        RECT 2.3500 2.0400 2.5400 2.0800 ;
        RECT 2.8700 2.0400 3.0600 2.0800 ;
        RECT 3.9150 2.0400 4.0850 2.0800 ;
        RECT 4.4750 2.0400 4.6450 2.0800 ;
        RECT 5.8500 1.8400 6.0600 2.0800 ;
        RECT 0.0750 1.7150 0.1750 2.0800 ;
        RECT 6.4250 1.5100 6.5250 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5000 1.4500 2.9500 1.5500 ;
    END
    ANTENNAGATEAREA 0.111 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.8600 4.1500 1.2800 ;
    END
    ANTENNAGATEAREA 0.111 ;
  END C

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2800 1.0500 3.6600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2589 ;
  END S0
  OBS
    LAYER M1 ;
      RECT 0.8050 1.6450 1.5200 1.7350 ;
      RECT 1.1950 0.9350 1.2850 1.6450 ;
      RECT 0.8050 0.8450 1.2850 0.9350 ;
      RECT 1.1950 0.7750 1.2850 0.8450 ;
      RECT 1.1950 0.6850 1.9800 0.7750 ;
      RECT 1.8900 0.5650 1.9800 0.6850 ;
      RECT 0.2800 1.8300 2.0400 1.9200 ;
      RECT 0.3350 0.6450 0.9450 0.7350 ;
      RECT 0.8550 0.5950 0.9450 0.6450 ;
      RECT 0.8550 0.5050 1.5200 0.5950 ;
      RECT 0.6050 0.7350 0.6950 1.8300 ;
      RECT 0.3350 0.7350 0.4350 0.9000 ;
      RECT 0.3350 0.4600 0.4350 0.6450 ;
      RECT 1.5550 1.2500 3.3350 1.3400 ;
      RECT 2.0800 1.4700 2.2900 1.5600 ;
      RECT 2.0800 1.3400 2.1700 1.4700 ;
      RECT 1.5550 1.0850 1.6450 1.2500 ;
      RECT 2.0800 0.8000 2.1700 1.2500 ;
      RECT 2.0800 0.4100 2.2300 0.8000 ;
      RECT 2.5950 1.6500 3.2600 1.7400 ;
      RECT 3.1700 1.5450 3.2600 1.6500 ;
      RECT 3.1700 1.4550 3.5350 1.5450 ;
      RECT 3.4450 1.3600 3.5350 1.4550 ;
      RECT 3.4450 1.2700 3.8400 1.3600 ;
      RECT 3.7500 0.9300 3.8400 1.2700 ;
      RECT 2.6600 0.8400 3.8400 0.9300 ;
      RECT 2.6600 0.4900 2.7500 0.8400 ;
      RECT 3.6450 1.4500 4.3900 1.5400 ;
      RECT 4.3000 0.7500 4.3900 1.4500 ;
      RECT 3.1000 0.6600 4.3900 0.7500 ;
      RECT 2.2400 1.8300 5.5100 1.9200 ;
      RECT 4.6600 0.9300 4.7500 1.8300 ;
      RECT 4.6600 0.8400 4.9500 0.9300 ;
      RECT 2.2400 1.7400 2.3300 1.8300 ;
      RECT 1.6300 1.6500 2.3300 1.7400 ;
      RECT 1.6300 1.5400 1.7200 1.6500 ;
      RECT 1.3750 1.4500 1.7200 1.5400 ;
      RECT 1.3750 0.9550 1.4650 1.4500 ;
      RECT 1.3750 0.8650 1.7800 0.9550 ;
      RECT 5.0600 0.8150 5.5100 0.9050 ;
      RECT 3.3700 1.6500 4.5700 1.7400 ;
      RECT 4.4800 0.7500 4.5700 1.6500 ;
      RECT 4.4800 0.6600 5.1500 0.7500 ;
      RECT 5.0600 0.7500 5.1500 0.8150 ;
      RECT 4.4800 0.5700 4.5700 0.6600 ;
      RECT 3.3650 0.4800 4.5700 0.5700 ;
      RECT 5.0600 0.9050 5.1500 1.0200 ;
      RECT 4.8400 1.0200 5.1500 1.1100 ;
      RECT 4.8400 1.1100 4.9300 1.7200 ;
      RECT 5.0250 1.4600 5.7800 1.5500 ;
      RECT 5.6900 0.9050 5.7800 1.4600 ;
      RECT 5.6100 0.7000 5.7800 0.9050 ;
      RECT 5.0250 1.2200 5.1150 1.4600 ;
      RECT 5.0550 1.6400 6.0650 1.7300 ;
      RECT 5.9750 0.5700 6.0650 1.6400 ;
      RECT 5.0400 0.4800 6.0650 0.5700 ;
  END
END MXT4_X1P4M_A12TH

MACRO MXT4_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9450 ;
        RECT 0.5650 0.3200 0.7550 0.5850 ;
        RECT 2.9450 0.3200 3.0450 0.7050 ;
        RECT 3.4600 0.3200 3.5600 0.5350 ;
        RECT 7.4350 0.3200 7.6250 0.3700 ;
        RECT 8.0200 0.3200 8.1200 0.6850 ;
    END
  END VSS

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6100 1.0500 7.1000 1.1500 ;
    END
    ANTENNAGATEAREA 0.1611 ;
  END S1

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 1.2500 0.5100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.2300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0500 0.9550 8.1500 1.2500 ;
        RECT 7.7650 1.2500 8.1500 1.3500 ;
        RECT 7.7650 0.8550 8.1500 0.9550 ;
        RECT 7.7650 1.3500 7.8650 1.7400 ;
        RECT 7.7650 0.5000 7.8650 0.8550 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 7.4700 1.8800 7.6400 2.0800 ;
        RECT 8.0200 1.7750 8.1200 2.0800 ;
        RECT 0.0750 1.7500 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0100 0.8500 3.5900 0.9500 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8600 5.1500 1.2800 ;
    END
    ANTENNAGATEAREA 0.1338 ;
  END C

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8300 1.0500 4.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.315 ;
  END S0
  OBS
    LAYER M1 ;
      RECT 0.3400 1.8300 2.2700 1.9200 ;
      RECT 2.1800 1.6750 2.2700 1.8300 ;
      RECT 0.6050 0.6850 1.8100 0.7750 ;
      RECT 0.6050 0.9500 0.6950 1.8300 ;
      RECT 0.3350 0.8600 0.6950 0.9500 ;
      RECT 0.6050 0.7750 0.6950 0.8600 ;
      RECT 0.3400 1.5200 0.4300 1.8300 ;
      RECT 0.3350 0.4950 0.4350 0.8600 ;
      RECT 0.8300 1.6450 1.8150 1.7350 ;
      RECT 1.1600 1.3550 1.2500 1.6450 ;
      RECT 1.1600 1.2650 1.4350 1.3550 ;
      RECT 1.3450 0.9550 1.4350 1.2650 ;
      RECT 0.8300 0.8650 2.2700 0.9550 ;
      RECT 2.1800 0.6800 2.2700 0.8650 ;
      RECT 1.7250 1.2550 3.9950 1.3450 ;
      RECT 2.6900 1.3450 2.7800 1.7100 ;
      RECT 2.6300 0.7450 2.7200 1.2550 ;
      RECT 2.6300 0.5150 2.7850 0.7450 ;
      RECT 3.2100 1.4500 4.3400 1.5400 ;
      RECT 4.2500 1.3600 4.3400 1.4500 ;
      RECT 4.2500 1.2700 4.7200 1.3600 ;
      RECT 4.6300 0.9300 4.7200 1.2700 ;
      RECT 3.7250 0.8400 4.7200 0.9300 ;
      RECT 3.7250 0.7500 3.8150 0.8400 ;
      RECT 3.2100 0.6600 3.8150 0.7500 ;
      RECT 3.2100 1.5400 3.3000 1.7400 ;
      RECT 3.2100 0.5100 3.3000 0.6600 ;
      RECT 4.4550 1.4500 5.4350 1.5400 ;
      RECT 5.3450 0.7500 5.4350 1.4500 ;
      RECT 3.9250 0.6600 5.4350 0.7500 ;
      RECT 2.4400 1.8300 6.8100 1.9200 ;
      RECT 6.7200 1.6400 6.8100 1.8300 ;
      RECT 5.7500 0.9300 5.8400 1.8300 ;
      RECT 5.7500 0.8400 6.3200 0.9300 ;
      RECT 2.4400 1.5550 2.5300 1.8300 ;
      RECT 1.3600 1.4650 2.5300 1.5550 ;
      RECT 1.5250 1.1500 1.6150 1.4650 ;
      RECT 1.5250 1.0600 2.5300 1.1500 ;
      RECT 2.4400 0.5700 2.5300 1.0600 ;
      RECT 1.3400 0.4800 2.5300 0.5700 ;
      RECT 5.5700 0.6600 6.8700 0.7500 ;
      RECT 3.6750 1.6500 5.6600 1.7400 ;
      RECT 5.5700 0.7500 5.6600 1.6500 ;
      RECT 6.4300 0.7500 6.5200 1.0200 ;
      RECT 5.5700 0.5700 5.6600 0.6600 ;
      RECT 6.1200 1.0200 6.5200 1.1100 ;
      RECT 3.6700 0.4800 5.6600 0.5700 ;
      RECT 6.1200 1.1100 6.2100 1.4500 ;
      RECT 6.1200 1.4500 6.3500 1.5400 ;
      RECT 7.2300 1.3550 7.3200 1.5050 ;
      RECT 6.3200 1.2650 7.3900 1.3550 ;
      RECT 7.3000 0.8850 7.3900 1.2650 ;
      RECT 7.1700 0.7950 7.3900 0.8850 ;
      RECT 6.3200 1.2200 6.4900 1.2650 ;
      RECT 7.5100 1.0600 7.8450 1.1600 ;
      RECT 6.4600 1.4550 7.0700 1.5450 ;
      RECT 6.9800 1.5450 7.0700 1.6300 ;
      RECT 6.9800 1.6300 7.6000 1.7200 ;
      RECT 7.5100 1.1600 7.6000 1.6300 ;
      RECT 7.5100 0.5700 7.6000 1.0600 ;
      RECT 5.8550 0.4800 7.6000 0.5700 ;
      RECT 5.9400 1.6500 6.5500 1.7400 ;
      RECT 6.4600 1.5450 6.5500 1.6500 ;
      RECT 5.9400 1.5250 6.0300 1.6500 ;
  END
END MXT4_X2M_A12TH

MACRO MXT4_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 0.0650 0.3200 0.1750 0.7150 ;
        RECT 0.5650 0.3200 0.7350 0.5100 ;
        RECT 1.1300 0.3200 1.2300 0.5150 ;
        RECT 2.7050 0.3200 2.8050 0.7200 ;
        RECT 3.2500 0.3200 3.3500 0.7500 ;
        RECT 3.7950 0.3200 3.8950 0.5650 ;
        RECT 7.7750 0.3200 7.9650 0.3700 ;
        RECT 8.3400 0.3200 8.4400 0.6850 ;
    END
  END VSS

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9500 1.0500 7.3850 1.1500 ;
    END
    ANTENNAGATEAREA 0.2181 ;
  END S1

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.4700 1.1500 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9400 1.0500 1.3900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0800 1.2500 8.7100 1.3500 ;
        RECT 8.0800 1.3500 8.1800 1.7400 ;
        RECT 8.6100 1.3500 8.7100 1.7400 ;
        RECT 8.6100 0.9550 8.7100 1.2500 ;
        RECT 8.0800 0.8550 8.7100 0.9550 ;
        RECT 8.0800 0.5300 8.1800 0.8550 ;
        RECT 8.6100 0.5300 8.7100 0.8550 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 7.7850 1.8800 7.9550 2.0800 ;
        RECT 8.3400 1.7750 8.4400 2.0800 ;
        RECT 0.0850 1.7500 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3700 1.0500 3.7900 1.1500 ;
        RECT 3.3700 1.1500 3.4700 1.3500 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 0.8600 5.5500 1.2800 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END C

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0500 3.2600 1.1500 ;
        RECT 3.1700 0.9600 3.2600 1.0500 ;
        RECT 3.1700 0.8700 3.9900 0.9600 ;
        RECT 3.9000 0.9600 3.9900 1.0250 ;
        RECT 3.9000 1.0250 5.1600 1.1150 ;
    END
    ANTENNAGATEAREA 0.4284 ;
  END S0
  OBS
    LAYER M1 ;
      RECT 0.8650 1.6450 1.8200 1.7350 ;
      RECT 0.8650 1.3900 0.9550 1.6450 ;
      RECT 0.7450 1.3000 0.9550 1.3900 ;
      RECT 0.7450 0.8400 2.2750 0.9300 ;
      RECT 2.1850 0.7200 2.2750 0.8400 ;
      RECT 0.7450 0.9300 0.8350 1.3000 ;
      RECT 0.5650 1.8300 2.3350 1.9200 ;
      RECT 0.3050 0.6600 1.8150 0.7500 ;
      RECT 0.3450 1.5750 0.4350 1.8950 ;
      RECT 0.3050 0.4450 0.4750 0.6600 ;
      RECT 0.5650 1.5750 0.6550 1.8300 ;
      RECT 0.3450 1.4850 0.6550 1.5750 ;
      RECT 0.5650 0.7500 0.6550 1.4850 ;
      RECT 3.5850 1.2600 4.4650 1.3500 ;
      RECT 4.0650 1.2100 4.4650 1.2600 ;
      RECT 1.7350 1.2300 1.9050 1.2600 ;
      RECT 2.6400 1.3500 2.7300 1.6250 ;
      RECT 1.7350 1.2600 2.7300 1.3500 ;
      RECT 2.6400 0.9300 2.7300 1.2600 ;
      RECT 2.6400 0.8400 3.0750 0.9300 ;
      RECT 2.9850 0.5050 3.0750 0.8400 ;
      RECT 3.2550 1.4500 3.6750 1.5400 ;
      RECT 3.5850 1.3500 3.6750 1.4500 ;
      RECT 2.6400 1.6250 3.3450 1.7150 ;
      RECT 3.2550 1.5400 3.3450 1.6250 ;
      RECT 3.8050 1.4500 4.6700 1.5400 ;
      RECT 4.5800 1.3200 4.6700 1.4500 ;
      RECT 4.5800 1.2300 5.3600 1.3200 ;
      RECT 5.2700 0.9300 5.3600 1.2300 ;
      RECT 4.0800 0.8400 5.3600 0.9300 ;
      RECT 4.0800 0.7800 4.1700 0.8400 ;
      RECT 3.4850 0.6900 4.1700 0.7800 ;
      RECT 3.4650 1.6500 3.8950 1.7400 ;
      RECT 3.8050 1.5400 3.8950 1.6500 ;
      RECT 3.4850 0.4750 3.6550 0.6900 ;
      RECT 4.7800 1.4400 5.7350 1.5300 ;
      RECT 5.6450 0.7500 5.7350 1.4400 ;
      RECT 4.2800 0.6600 5.7350 0.7500 ;
      RECT 5.8250 0.6600 7.1550 0.7500 ;
      RECT 4.0050 1.6500 5.9150 1.7400 ;
      RECT 5.8250 0.7500 5.9150 1.6500 ;
      RECT 6.7500 0.7500 6.8400 1.0400 ;
      RECT 5.8250 0.5700 5.9150 0.6600 ;
      RECT 6.2450 1.0400 6.8400 1.1300 ;
      RECT 3.9900 0.4800 5.9150 0.5700 ;
      RECT 6.2450 1.1300 6.3350 1.4250 ;
      RECT 6.2450 1.4250 6.6350 1.5150 ;
      RECT 2.4450 1.8300 7.4050 1.9200 ;
      RECT 6.0050 0.9300 6.0950 1.8300 ;
      RECT 6.0050 0.8400 6.6350 0.9300 ;
      RECT 2.4450 1.5550 2.5350 1.8300 ;
      RECT 1.3450 1.4650 2.5350 1.5550 ;
      RECT 1.5100 1.1400 1.6100 1.4650 ;
      RECT 1.5100 1.0400 2.5500 1.1400 ;
      RECT 2.4500 0.5700 2.5500 1.0400 ;
      RECT 1.3400 0.4800 2.5500 0.5700 ;
      RECT 6.7550 1.4150 7.6350 1.5050 ;
      RECT 7.5450 0.7200 7.6350 1.4150 ;
      RECT 6.7550 1.3200 6.8450 1.4150 ;
      RECT 6.5750 1.2300 6.8450 1.3200 ;
      RECT 7.8250 1.0500 8.4550 1.1500 ;
      RECT 6.1850 1.6300 7.9150 1.7200 ;
      RECT 7.8250 1.1500 7.9150 1.6300 ;
      RECT 7.8250 0.5700 7.9150 1.0500 ;
      RECT 6.1600 0.4800 7.9150 0.5700 ;
      RECT 7.2650 0.5700 7.3550 0.9050 ;
  END
END MXT4_X3M_A12TH

MACRO M2SDFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.4050 0.3200 0.5050 0.7100 ;
        RECT 2.6500 0.3200 2.8200 0.4700 ;
        RECT 3.1500 0.3200 3.3200 0.4800 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0774 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7250 1.0500 3.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5350 1.4500 2.9550 1.5500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 0.8200 7.3700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.7800 6.5500 1.3150 ;
        RECT 6.4500 1.3150 6.6350 1.4150 ;
        RECT 6.4500 0.6900 6.6700 0.7800 ;
        RECT 6.5350 1.4150 6.6350 1.7250 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 2.6400 1.8450 2.8100 2.0800 ;
        RECT 0.3300 1.7550 0.5000 2.0800 ;
        RECT 3.1800 1.5600 3.2900 2.0800 ;
        RECT 1.6300 1.4200 1.7300 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8650 1.5800 1.2550 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 3.6750 1.5000 3.9200 1.5900 ;
      RECT 3.8300 0.7700 3.9200 1.5000 ;
      RECT 3.8300 0.6800 4.5900 0.7700 ;
      RECT 4.5000 0.7700 4.5900 0.9750 ;
      RECT 4.4550 0.9750 4.5900 1.1200 ;
      RECT 4.4550 1.1200 4.5450 1.3650 ;
      RECT 4.1250 1.4850 4.7700 1.5750 ;
      RECT 4.1250 1.1650 4.2150 1.4850 ;
      RECT 4.6800 0.7700 4.7700 1.4850 ;
      RECT 4.6800 0.6800 4.8500 0.7700 ;
      RECT 4.8550 1.6400 5.4150 1.7300 ;
      RECT 5.3250 0.7700 5.4150 1.6400 ;
      RECT 5.1200 0.6800 5.8350 0.7700 ;
      RECT 5.7450 0.7700 5.8350 0.9850 ;
      RECT 5.7450 0.9850 5.9550 1.0750 ;
      RECT 5.8650 1.0750 5.9550 1.4250 ;
      RECT 5.5250 1.6400 6.3350 1.7300 ;
      RECT 5.5250 1.2750 5.6150 1.6400 ;
      RECT 6.2450 0.7550 6.3350 1.6400 ;
      RECT 5.9650 0.6650 6.3350 0.7550 ;
      RECT 3.6500 0.4800 6.8800 0.5700 ;
      RECT 6.7900 0.5700 6.8800 1.6100 ;
      RECT 5.1150 1.0400 5.2050 1.5300 ;
      RECT 4.9400 0.9500 5.2050 1.0400 ;
      RECT 4.9400 0.5700 5.0300 0.9500 ;
      RECT 3.6500 0.5700 3.7400 1.3850 ;
      RECT 3.9250 0.4100 4.0950 0.4800 ;
      RECT 6.9700 1.5000 7.5550 1.5900 ;
      RECT 6.9700 0.6100 7.5550 0.7000 ;
      RECT 3.7850 1.8300 7.0600 1.9200 ;
      RECT 6.9700 1.5900 7.0600 1.8300 ;
      RECT 6.9700 0.7000 7.0600 1.5000 ;
      RECT 4.7950 1.9200 4.9650 1.9650 ;
      RECT 0.7000 1.3750 0.9400 1.4650 ;
      RECT 0.8400 0.6650 0.9400 1.3750 ;
      RECT 0.7050 0.5750 0.9400 0.6650 ;
      RECT 0.7850 1.8800 1.1200 1.9700 ;
      RECT 0.7850 1.6450 0.8750 1.8800 ;
      RECT 0.4400 1.5550 0.8750 1.6450 ;
      RECT 0.4400 1.5450 0.5300 1.5550 ;
      RECT 0.0500 1.4550 0.5300 1.5450 ;
      RECT 0.0500 1.5450 0.1700 1.8900 ;
      RECT 0.0500 0.6550 0.1400 1.4550 ;
      RECT 0.0500 0.5650 0.2400 0.6550 ;
      RECT 1.3350 1.4400 1.4250 1.7800 ;
      RECT 1.2250 1.3500 1.4250 1.4400 ;
      RECT 1.2250 0.7500 1.3150 1.3500 ;
      RECT 1.2250 0.6600 1.4400 0.7500 ;
      RECT 1.8850 1.3050 1.9750 1.9800 ;
      RECT 1.7950 1.2150 1.9750 1.3050 ;
      RECT 1.7950 0.5700 1.8850 1.2150 ;
      RECT 1.0300 0.4800 1.8850 0.5700 ;
      RECT 1.0300 0.5700 1.1200 1.7750 ;
      RECT 2.9400 1.7450 3.0300 1.9300 ;
      RECT 2.3250 1.6550 3.0300 1.7450 ;
      RECT 2.3250 0.7800 3.1500 0.8700 ;
      RECT 2.3250 0.8700 2.4150 1.6550 ;
      RECT 2.1450 0.5800 3.3500 0.6700 ;
      RECT 3.2600 0.6700 3.3500 1.3250 ;
      RECT 2.1450 0.6700 2.2350 1.9800 ;
      RECT 3.4500 0.4250 3.5400 1.7550 ;
  END
END M2SDFFQN_X1M_A12TH

MACRO M2SDFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6800 ;
        RECT 2.6150 0.3200 2.7850 0.5050 ;
        RECT 3.2400 0.3200 3.4100 0.4800 ;
        RECT 7.3300 0.3200 7.5000 0.5000 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.1002 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7550 1.4500 3.2050 1.5500 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0500 2.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.8350 7.5550 1.2600 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.8100 6.7500 1.2500 ;
        RECT 6.5100 1.2500 6.7500 1.3500 ;
        RECT 6.4500 0.7100 6.7500 0.8100 ;
        RECT 6.5150 1.3500 6.6050 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 0.3150 1.8750 0.4850 2.0800 ;
        RECT 2.5900 1.8650 2.7600 2.0800 ;
        RECT 3.2550 1.7200 3.3650 2.0800 ;
        RECT 1.5350 1.5500 1.6350 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 6.0650 1.0700 6.5400 1.1600 ;
      RECT 6.0050 1.3900 6.0950 1.6900 ;
      RECT 5.6050 1.3000 6.1550 1.3900 ;
      RECT 6.0650 1.1600 6.1550 1.3000 ;
      RECT 5.6050 1.0400 5.6950 1.3000 ;
      RECT 6.0650 0.9300 6.1550 1.0700 ;
      RECT 5.9650 0.8400 6.1550 0.9300 ;
      RECT 3.7250 0.4800 7.1150 0.5700 ;
      RECT 7.0250 0.5700 7.1150 1.5300 ;
      RECT 5.2250 1.0500 5.3150 1.5050 ;
      RECT 4.9300 0.9600 5.3150 1.0500 ;
      RECT 4.9300 0.5700 5.0200 0.9600 ;
      RECT 3.7250 0.5700 3.8150 1.4050 ;
      RECT 3.9700 0.4250 4.1400 0.4800 ;
      RECT 7.0100 1.6450 7.7200 1.7350 ;
      RECT 7.6300 1.5250 7.7200 1.6450 ;
      RECT 7.2150 0.6100 7.7200 0.7000 ;
      RECT 7.6300 0.4450 7.7200 0.6100 ;
      RECT 3.9850 1.8300 7.1000 1.9200 ;
      RECT 7.0100 1.7350 7.1000 1.8300 ;
      RECT 7.2150 0.7000 7.3050 1.6450 ;
      RECT 4.9000 1.4950 4.9900 1.8300 ;
      RECT 4.9000 1.3250 5.0400 1.4950 ;
      RECT 0.5900 1.3200 0.7300 1.5100 ;
      RECT 0.6400 0.6900 0.7300 1.3200 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0950 1.6200 0.9100 1.7100 ;
      RECT 0.8200 1.0600 0.9100 1.6200 ;
      RECT 0.2550 0.8700 0.3450 1.6200 ;
      RECT 0.0950 0.7800 0.3450 0.8700 ;
      RECT 0.0950 1.7100 0.1850 1.9900 ;
      RECT 0.0950 0.4800 0.1850 0.7800 ;
      RECT 1.2600 0.7550 1.3500 1.9050 ;
      RECT 1.1550 0.6650 1.3500 0.7550 ;
      RECT 0.8900 0.4800 1.9000 0.5700 ;
      RECT 1.8100 0.5700 1.9000 1.9150 ;
      RECT 1.0000 0.9150 1.0900 1.8850 ;
      RECT 0.8900 0.8250 1.0900 0.9150 ;
      RECT 0.8900 0.5700 0.9800 0.8250 ;
      RECT 2.9100 1.7600 3.0000 1.9800 ;
      RECT 2.2500 1.6700 3.0000 1.7600 ;
      RECT 2.2500 0.8250 3.1650 0.9150 ;
      RECT 2.2500 0.9150 2.3400 1.6700 ;
      RECT 2.0700 0.6250 3.4250 0.7150 ;
      RECT 3.3350 0.7150 3.4250 1.3450 ;
      RECT 2.0700 0.7150 2.1600 1.9150 ;
      RECT 2.0700 0.5200 2.1600 0.6250 ;
      RECT 3.5400 0.4650 3.6300 1.8300 ;
      RECT 3.8000 1.6200 3.8900 1.9250 ;
      RECT 3.8000 1.5300 3.9950 1.6200 ;
      RECT 3.9050 0.7550 3.9950 1.5300 ;
      RECT 3.9050 0.6650 4.6100 0.7550 ;
      RECT 4.5200 0.7550 4.6100 1.1750 ;
      RECT 4.2100 1.5700 4.8100 1.6600 ;
      RECT 4.2100 1.1150 4.3000 1.5700 ;
      RECT 4.7200 0.6650 4.8100 1.5700 ;
      RECT 5.0800 1.6300 5.5150 1.7200 ;
      RECT 5.4250 0.7550 5.5150 1.6300 ;
      RECT 5.1200 0.6650 5.8750 0.7550 ;
      RECT 5.1200 0.7550 5.2100 0.8350 ;
      RECT 5.7850 0.7550 5.8750 1.0900 ;
      RECT 5.7850 1.0900 5.9750 1.1800 ;
  END
END M2SDFFQN_X2M_A12TH

MACRO M2SDFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.0450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6800 ;
        RECT 2.6150 0.3200 2.7850 0.5250 ;
        RECT 3.2400 0.3200 3.4100 0.5300 ;
        RECT 4.4200 0.3200 4.5900 0.3900 ;
        RECT 7.5300 0.3200 7.7000 0.5200 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.1002 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7550 1.4500 3.2050 1.5500 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0500 2.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8350 0.8350 7.9500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8500 0.8150 6.9500 1.2500 ;
        RECT 6.5100 1.2500 7.1250 1.3500 ;
        RECT 6.4500 0.7150 7.1600 0.8150 ;
        RECT 6.5100 1.3500 6.6000 1.7200 ;
        RECT 7.0250 1.3500 7.1250 1.7250 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.0450 2.7200 ;
        RECT 0.3150 1.8750 0.4850 2.0800 ;
        RECT 2.5850 1.8500 2.7550 2.0800 ;
        RECT 7.5050 1.7750 7.6750 2.0800 ;
        RECT 3.2550 1.6350 3.3650 2.0800 ;
        RECT 1.5350 1.5700 1.6350 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 2.0700 0.6250 3.4250 0.7150 ;
      RECT 3.3350 0.7150 3.4250 1.3450 ;
      RECT 2.0700 0.7150 2.1600 1.8550 ;
      RECT 2.0700 0.5200 2.1600 0.6250 ;
      RECT 3.5400 0.4650 3.6300 1.9000 ;
      RECT 3.8000 1.6200 3.8900 1.9400 ;
      RECT 3.8000 1.5300 3.9950 1.6200 ;
      RECT 3.9050 0.7550 3.9950 1.5300 ;
      RECT 3.9050 0.6650 4.6100 0.7550 ;
      RECT 4.5200 0.7550 4.6100 1.1750 ;
      RECT 4.2100 1.5700 4.8100 1.6600 ;
      RECT 4.2100 1.1150 4.3000 1.5700 ;
      RECT 4.7200 0.6650 4.8100 1.5700 ;
      RECT 5.0800 1.6300 5.4950 1.7200 ;
      RECT 5.4050 1.1800 5.4950 1.6300 ;
      RECT 5.4050 1.0900 5.9100 1.1800 ;
      RECT 5.4050 0.7550 5.4950 1.0900 ;
      RECT 5.1200 0.6650 5.5150 0.7550 ;
      RECT 5.1200 0.7550 5.2100 0.8350 ;
      RECT 6.0000 1.0700 6.7400 1.1600 ;
      RECT 5.5850 1.6150 6.0900 1.7050 ;
      RECT 5.5850 1.3200 5.6750 1.6150 ;
      RECT 6.0000 1.1600 6.0900 1.6150 ;
      RECT 6.0000 0.7500 6.0900 1.0700 ;
      RECT 3.7250 0.4800 7.3700 0.5700 ;
      RECT 7.2800 0.5700 7.3700 1.5000 ;
      RECT 5.2250 1.0500 5.3150 1.5050 ;
      RECT 4.9200 0.9600 5.3150 1.0500 ;
      RECT 4.9200 0.5700 5.0100 0.9600 ;
      RECT 3.7250 0.5700 3.8150 1.4050 ;
      RECT 3.9700 0.4250 4.1400 0.4800 ;
      RECT 7.2650 1.5900 7.9200 1.6800 ;
      RECT 7.8300 1.4950 7.9200 1.5900 ;
      RECT 7.4800 0.6100 7.9200 0.7000 ;
      RECT 7.8300 0.4450 7.9200 0.6100 ;
      RECT 7.4800 0.7000 7.5700 1.5900 ;
      RECT 3.9850 1.8300 7.3550 1.9200 ;
      RECT 7.2650 1.6800 7.3550 1.8300 ;
      RECT 4.9000 1.4950 4.9900 1.8300 ;
      RECT 4.9000 1.3250 5.0400 1.4950 ;
      RECT 0.5900 1.3200 0.7300 1.5150 ;
      RECT 0.6400 0.6900 0.7300 1.3200 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0950 1.5600 0.4800 1.6500 ;
      RECT 0.3900 1.6500 0.4800 1.6750 ;
      RECT 0.3900 1.6750 0.9100 1.7650 ;
      RECT 0.8200 1.0350 0.9100 1.6750 ;
      RECT 0.2550 0.8750 0.3450 1.5600 ;
      RECT 0.0950 0.7850 0.3450 0.8750 ;
      RECT 0.0950 1.6500 0.1850 1.9800 ;
      RECT 0.0950 0.4850 0.1850 0.7850 ;
      RECT 1.2600 0.7550 1.3500 1.8650 ;
      RECT 1.1550 0.6650 1.3500 0.7550 ;
      RECT 0.8900 0.4800 1.9000 0.5700 ;
      RECT 1.8100 0.5700 1.9000 1.8550 ;
      RECT 1.0000 0.9150 1.0900 1.8450 ;
      RECT 0.8900 0.8250 1.0900 0.9150 ;
      RECT 0.8900 0.5700 0.9800 0.8250 ;
      RECT 2.9300 1.7450 3.0200 1.9900 ;
      RECT 2.2500 1.6550 3.0200 1.7450 ;
      RECT 2.2500 0.8250 3.1650 0.9150 ;
      RECT 2.2500 0.9150 2.3400 1.6550 ;
  END
END M2SDFFQN_X3M_A12TH

MACRO M2SDFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.3350 0.3200 0.5050 0.6700 ;
        RECT 2.6250 0.3200 2.7950 0.4850 ;
        RECT 3.0650 0.3200 3.1750 0.4500 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8400 0.5950 1.3600 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8100 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5800 1.0500 3.0000 1.1500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SE

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8450 1.5500 1.2650 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D0

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2400 0.8350 7.3550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.8650 6.5500 1.4500 ;
        RECT 6.4500 1.4500 6.6400 1.5500 ;
        RECT 6.4500 0.7650 6.6750 0.8650 ;
        RECT 6.5400 1.5500 6.6400 1.6950 ;
    END
    ANTENNADIFFAREA 0.1224 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 2.5800 1.8500 2.7500 2.0800 ;
        RECT 0.3950 1.7000 0.4950 2.0800 ;
        RECT 3.1550 1.5050 3.2750 2.0800 ;
        RECT 1.5550 1.4950 1.6550 2.0800 ;
    END
  END VDD

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.4500 2.8700 1.5500 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SI
  OBS
    LAYER M1 ;
      RECT 4.8700 1.5550 5.3450 1.6450 ;
      RECT 5.2550 0.7700 5.3450 1.5550 ;
      RECT 5.1100 0.6800 6.3550 0.7700 ;
      RECT 5.7400 0.7700 5.8300 1.1100 ;
      RECT 6.2650 0.7700 6.3550 1.2450 ;
      RECT 5.7400 1.1100 5.9600 1.2000 ;
      RECT 5.8700 1.2000 5.9600 1.3200 ;
      RECT 3.6350 0.4800 6.8650 0.5700 ;
      RECT 6.7750 0.5700 6.8650 1.6550 ;
      RECT 4.9300 1.3000 5.1350 1.3900 ;
      RECT 4.9300 0.5700 5.0200 1.3000 ;
      RECT 3.6350 0.5700 3.7250 1.4350 ;
      RECT 3.8900 0.4350 4.0600 0.4800 ;
      RECT 6.9600 1.5000 7.5200 1.5900 ;
      RECT 7.4300 1.5900 7.5200 1.6900 ;
      RECT 6.9600 0.6100 7.5200 0.7000 ;
      RECT 7.4300 0.5100 7.5200 0.6100 ;
      RECT 3.8050 1.8200 7.0500 1.9100 ;
      RECT 6.9600 1.5900 7.0500 1.8200 ;
      RECT 6.9600 0.7000 7.0500 1.5000 ;
      RECT 0.7800 0.7300 0.8800 1.7150 ;
      RECT 0.6350 0.6400 0.8800 0.7300 ;
      RECT 0.8750 1.9150 1.0850 1.9650 ;
      RECT 0.5950 1.8250 1.0850 1.9150 ;
      RECT 0.5950 1.5900 0.6850 1.8250 ;
      RECT 0.0500 1.5000 0.6850 1.5900 ;
      RECT 0.0500 1.5900 0.1700 1.7300 ;
      RECT 0.0500 0.7300 0.1400 1.5000 ;
      RECT 0.0500 0.5600 0.2000 0.7300 ;
      RECT 1.3000 1.4850 1.3900 1.7000 ;
      RECT 1.1850 1.3950 1.3900 1.4850 ;
      RECT 1.1850 0.7500 1.2750 1.3950 ;
      RECT 1.1850 0.6600 1.3600 0.7500 ;
      RECT 0.9700 0.4800 1.9000 0.5700 ;
      RECT 1.8100 0.5700 1.9000 1.9150 ;
      RECT 0.9700 1.6050 1.1900 1.6950 ;
      RECT 0.9700 0.5700 1.0600 1.6050 ;
      RECT 2.8950 1.7500 2.9850 1.9600 ;
      RECT 2.2500 1.6600 2.9850 1.7500 ;
      RECT 2.2500 0.8600 3.0850 0.9500 ;
      RECT 2.9950 0.7600 3.0850 0.8600 ;
      RECT 2.2500 0.9500 2.3400 1.6600 ;
      RECT 2.0700 0.5750 3.3400 0.6650 ;
      RECT 3.2500 0.6650 3.3400 1.3600 ;
      RECT 2.0700 0.6650 2.1600 1.9150 ;
      RECT 3.4500 0.6050 3.5400 1.6950 ;
      RECT 3.6900 1.5550 3.9050 1.6450 ;
      RECT 3.8150 0.7700 3.9050 1.5550 ;
      RECT 3.8150 0.6800 4.5800 0.7700 ;
      RECT 4.4900 0.7700 4.5800 1.2950 ;
      RECT 4.1500 1.5250 4.7600 1.6150 ;
      RECT 4.1500 1.1100 4.2400 1.5250 ;
      RECT 4.6700 0.7700 4.7600 1.5250 ;
      RECT 4.6700 0.6800 4.8400 0.7700 ;
      RECT 5.4950 1.5250 6.1750 1.6150 ;
      RECT 5.4950 0.9650 5.5850 1.5250 ;
      RECT 6.0850 0.9550 6.1750 1.5250 ;
      RECT 5.9750 0.8650 6.1750 0.9550 ;
  END
END M2SDFFQ_X0P5M_A12TH

MACRO M2SDFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.4050 0.3200 0.5050 0.7100 ;
        RECT 2.6500 0.3200 2.8200 0.4700 ;
        RECT 3.1900 0.3200 3.2800 0.4350 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0804 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7250 1.0500 3.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5350 1.4500 2.9550 1.5500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 0.8200 7.3700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.7550 6.5500 1.3150 ;
        RECT 6.4500 1.3150 6.6350 1.4150 ;
        RECT 6.4500 0.6650 6.6700 0.7550 ;
        RECT 6.5350 1.4150 6.6350 1.7200 ;
    END
    ANTENNADIFFAREA 0.2448 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 7.0700 2.0200 7.2400 2.0800 ;
        RECT 2.6400 1.8750 2.8100 2.0800 ;
        RECT 0.3700 1.7550 0.5400 2.0800 ;
        RECT 3.1800 1.5500 3.2900 2.0800 ;
        RECT 1.6300 1.4300 1.7300 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8650 1.5800 1.2550 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 3.6750 1.5000 3.9200 1.5900 ;
      RECT 3.8300 0.7700 3.9200 1.5000 ;
      RECT 3.8300 0.6800 4.5650 0.7700 ;
      RECT 4.4750 0.7700 4.5650 1.2750 ;
      RECT 4.1250 1.4700 4.7650 1.5600 ;
      RECT 4.1250 1.1650 4.2150 1.4700 ;
      RECT 4.6750 0.7700 4.7650 1.4700 ;
      RECT 4.6750 0.6800 4.8500 0.7700 ;
      RECT 5.5250 1.6400 6.1650 1.7300 ;
      RECT 5.5250 1.0850 5.6150 1.6400 ;
      RECT 6.0750 0.9500 6.1650 1.6400 ;
      RECT 5.9900 0.8600 6.1650 0.9500 ;
      RECT 4.8700 1.6400 5.4150 1.7300 ;
      RECT 5.3250 0.7700 5.4150 1.6400 ;
      RECT 5.1200 0.6800 6.3600 0.7700 ;
      RECT 5.7900 0.7700 5.8800 1.2950 ;
      RECT 6.2700 0.7700 6.3600 1.1600 ;
      RECT 3.6500 0.4800 6.8800 0.5700 ;
      RECT 6.7900 0.5700 6.8800 1.6100 ;
      RECT 5.1150 1.0350 5.2050 1.5300 ;
      RECT 4.9400 0.9450 5.2050 1.0350 ;
      RECT 4.9400 0.5700 5.0300 0.9450 ;
      RECT 3.6500 0.5700 3.7400 1.3850 ;
      RECT 3.9250 0.4100 4.0950 0.4800 ;
      RECT 6.9700 1.4800 7.5550 1.5700 ;
      RECT 6.9700 0.6300 7.5550 0.7200 ;
      RECT 3.7850 1.8300 7.0600 1.9200 ;
      RECT 6.9700 1.5700 7.0600 1.8300 ;
      RECT 6.9700 0.7200 7.0600 1.4800 ;
      RECT 4.7950 1.9200 4.9650 1.9650 ;
      RECT 0.7050 1.3750 0.9400 1.4650 ;
      RECT 0.8400 0.6650 0.9400 1.3750 ;
      RECT 0.7050 0.5750 0.9400 0.6650 ;
      RECT 0.7850 1.8800 1.1200 1.9700 ;
      RECT 0.7850 1.6450 0.8750 1.8800 ;
      RECT 0.4400 1.5550 0.8750 1.6450 ;
      RECT 0.4400 1.5450 0.5300 1.5550 ;
      RECT 0.0500 1.4550 0.5300 1.5450 ;
      RECT 0.0500 1.5450 0.1700 1.8700 ;
      RECT 0.0500 0.6550 0.1400 1.4550 ;
      RECT 0.0500 0.5650 0.2350 0.6550 ;
      RECT 1.3350 1.4550 1.4250 1.7800 ;
      RECT 1.2250 1.3650 1.4250 1.4550 ;
      RECT 1.2250 0.7500 1.3150 1.3650 ;
      RECT 1.2250 0.6600 1.4400 0.7500 ;
      RECT 1.8850 1.3550 1.9750 1.9600 ;
      RECT 1.7900 1.2650 1.9750 1.3550 ;
      RECT 1.7900 0.8650 1.8800 1.2650 ;
      RECT 1.7900 0.6950 1.8850 0.8650 ;
      RECT 1.7900 0.5700 1.8800 0.6950 ;
      RECT 1.0300 0.4800 1.8800 0.5700 ;
      RECT 1.0300 0.5700 1.1200 1.7750 ;
      RECT 2.9400 1.7600 3.0300 1.9600 ;
      RECT 2.3250 1.6700 3.0300 1.7600 ;
      RECT 2.3250 0.7800 3.1500 0.8700 ;
      RECT 2.3250 0.8700 2.4150 1.6700 ;
      RECT 2.1450 0.5800 3.3500 0.6700 ;
      RECT 3.2600 0.6700 3.3500 1.3250 ;
      RECT 2.1450 0.6700 2.2350 1.9700 ;
      RECT 3.4500 0.4250 3.5400 1.6650 ;
  END
END M2SDFFQ_X1M_A12TH

MACRO M2SDFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6800 ;
        RECT 2.6150 0.3200 2.7850 0.5050 ;
        RECT 3.2400 0.3200 3.4100 0.4800 ;
        RECT 7.3300 0.3200 7.5000 0.5000 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.5100 ;
    END
    ANTENNAGATEAREA 0.0864 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7550 1.4500 3.2050 1.5500 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0500 2.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.8350 7.5550 1.2600 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.8100 6.7500 1.2500 ;
        RECT 6.5100 1.2500 6.7500 1.3500 ;
        RECT 6.4500 0.7100 6.7500 0.8100 ;
        RECT 6.5100 1.3500 6.6000 1.7200 ;
    END
    ANTENNADIFFAREA 0.306 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 0.3150 1.8750 0.4850 2.0800 ;
        RECT 2.5900 1.8650 2.7600 2.0800 ;
        RECT 3.2550 1.7200 3.3650 2.0800 ;
        RECT 1.5350 1.5500 1.6350 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 6.2500 1.0700 6.5400 1.1600 ;
      RECT 5.0800 1.6300 5.5150 1.7200 ;
      RECT 5.4250 1.2050 5.5150 1.6300 ;
      RECT 5.4250 1.1150 5.9200 1.2050 ;
      RECT 5.4250 0.7700 5.5150 1.1150 ;
      RECT 5.4250 0.7550 6.3400 0.7700 ;
      RECT 6.2500 0.7700 6.3400 1.0700 ;
      RECT 5.1200 0.6800 6.3400 0.7550 ;
      RECT 5.1200 0.7550 5.2100 0.8350 ;
      RECT 5.1200 0.6650 5.5150 0.6800 ;
      RECT 3.7250 0.4800 7.1100 0.5700 ;
      RECT 7.0200 0.5700 7.1100 1.5300 ;
      RECT 5.2250 1.0500 5.3150 1.5050 ;
      RECT 4.9200 0.9600 5.3150 1.0500 ;
      RECT 4.9200 0.5700 5.0100 0.9600 ;
      RECT 3.7250 0.5700 3.8150 1.4050 ;
      RECT 3.9700 0.4250 4.1400 0.4800 ;
      RECT 7.0050 1.6450 7.7200 1.7350 ;
      RECT 7.6300 1.5250 7.7200 1.6450 ;
      RECT 7.2100 0.6100 7.7200 0.7000 ;
      RECT 7.6300 0.4450 7.7200 0.6100 ;
      RECT 3.9850 1.8300 7.0950 1.9200 ;
      RECT 7.0050 1.7350 7.0950 1.8300 ;
      RECT 7.2100 0.7000 7.3000 1.6450 ;
      RECT 4.9000 1.4950 4.9900 1.8300 ;
      RECT 4.9000 1.3250 5.0400 1.4950 ;
      RECT 0.5900 1.3200 0.7300 1.5150 ;
      RECT 0.6400 0.6900 0.7300 1.3200 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0550 1.6850 0.9100 1.7750 ;
      RECT 0.8200 1.0350 0.9100 1.6850 ;
      RECT 0.2550 0.8750 0.3450 1.6850 ;
      RECT 0.0950 0.7850 0.3450 0.8750 ;
      RECT 0.0950 0.4850 0.1850 0.7850 ;
      RECT 1.2600 0.7550 1.3500 1.8650 ;
      RECT 1.1550 0.6650 1.3500 0.7550 ;
      RECT 1.8100 1.4950 1.9450 1.8850 ;
      RECT 1.8550 0.6750 1.9450 1.4950 ;
      RECT 1.8100 0.5700 1.9450 0.6750 ;
      RECT 0.8900 0.4800 1.9450 0.5700 ;
      RECT 0.8900 0.5700 0.9800 0.8250 ;
      RECT 0.8900 0.8250 1.0900 0.9150 ;
      RECT 1.0000 0.9150 1.0900 1.8450 ;
      RECT 2.9100 1.7600 3.0000 1.9800 ;
      RECT 2.2500 1.6700 3.0000 1.7600 ;
      RECT 2.2500 0.8250 3.1650 0.9150 ;
      RECT 2.2500 0.9150 2.3400 1.6700 ;
      RECT 2.0700 0.6250 3.4250 0.7150 ;
      RECT 3.3350 0.7150 3.4250 1.3450 ;
      RECT 2.0700 0.7150 2.1600 1.8850 ;
      RECT 2.0700 0.5200 2.1600 0.6250 ;
      RECT 3.5400 0.4650 3.6300 1.8700 ;
      RECT 3.8000 1.6200 3.8900 1.9250 ;
      RECT 3.8000 1.5300 3.9950 1.6200 ;
      RECT 3.9050 0.7550 3.9950 1.5300 ;
      RECT 3.9050 0.6650 4.6100 0.7550 ;
      RECT 4.5200 0.7550 4.6100 1.1750 ;
      RECT 4.2100 1.5700 4.8100 1.6600 ;
      RECT 4.2100 1.1150 4.3000 1.5700 ;
      RECT 4.7200 0.6650 4.8100 1.5700 ;
      RECT 5.6050 1.6150 6.1550 1.7050 ;
      RECT 5.6050 1.3200 5.6950 1.6150 ;
      RECT 6.0650 0.9550 6.1550 1.6150 ;
      RECT 5.9450 0.8650 6.1550 0.9550 ;
  END
END M2SDFFQ_X2M_A12TH

MACRO M2SDFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.0450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6800 ;
        RECT 2.6150 0.3200 2.7850 0.5050 ;
        RECT 3.2400 0.3200 3.4100 0.5300 ;
        RECT 4.4100 0.3200 4.5800 0.3700 ;
        RECT 7.5300 0.3200 7.7000 0.4600 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.5050 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7550 1.4500 3.2050 1.5500 ;
    END
    ANTENNAGATEAREA 0.0621 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0500 2.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8350 0.8350 7.9500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8500 0.8150 6.9500 1.2500 ;
        RECT 6.5100 1.2500 7.1250 1.3500 ;
        RECT 6.4500 0.7150 7.1600 0.8150 ;
        RECT 6.5100 1.3500 6.6000 1.7200 ;
        RECT 7.0250 1.3500 7.1250 1.7250 ;
    END
    ANTENNADIFFAREA 0.6048 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.0450 2.7200 ;
        RECT 0.3150 1.8750 0.4850 2.0800 ;
        RECT 2.5900 1.8650 2.7600 2.0800 ;
        RECT 7.5050 1.8500 7.6750 2.0800 ;
        RECT 3.2550 1.6350 3.3650 2.0800 ;
        RECT 1.5350 1.5500 1.6350 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 2.0700 0.6250 3.4250 0.7150 ;
      RECT 3.3350 0.7150 3.4250 1.3450 ;
      RECT 2.0700 0.7150 2.1600 1.8850 ;
      RECT 2.0700 0.5200 2.1600 0.6250 ;
      RECT 3.5400 0.4650 3.6300 1.9000 ;
      RECT 3.8000 1.6200 3.8900 1.9400 ;
      RECT 3.8000 1.5300 3.9950 1.6200 ;
      RECT 3.9050 0.7550 3.9950 1.5300 ;
      RECT 3.9050 0.6650 4.6100 0.7550 ;
      RECT 4.5200 0.7550 4.6100 1.1750 ;
      RECT 4.2100 1.5700 4.8100 1.6600 ;
      RECT 4.2100 1.1150 4.3000 1.5700 ;
      RECT 4.7200 0.6650 4.8100 1.5700 ;
      RECT 5.6050 1.6150 6.1550 1.7050 ;
      RECT 5.6050 1.3200 5.6950 1.6150 ;
      RECT 6.0650 0.9550 6.1550 1.6150 ;
      RECT 5.9450 0.8650 6.1550 0.9550 ;
      RECT 6.2500 1.0700 6.7150 1.1600 ;
      RECT 5.0800 1.6300 5.5150 1.7200 ;
      RECT 5.4250 1.2050 5.5150 1.6300 ;
      RECT 5.4250 1.1150 5.9200 1.2050 ;
      RECT 5.4250 0.7700 5.5150 1.1150 ;
      RECT 5.4250 0.7550 6.3400 0.7700 ;
      RECT 6.2500 0.7700 6.3400 1.0700 ;
      RECT 5.1200 0.6800 6.3400 0.7550 ;
      RECT 5.1200 0.7550 5.2100 0.8350 ;
      RECT 5.1200 0.6650 5.5150 0.6800 ;
      RECT 3.7250 0.4800 7.3700 0.5700 ;
      RECT 7.2800 0.5700 7.3700 1.5300 ;
      RECT 5.2250 1.0500 5.3150 1.5050 ;
      RECT 4.9200 0.9600 5.3150 1.0500 ;
      RECT 4.9200 0.5700 5.0100 0.9600 ;
      RECT 3.7250 0.5700 3.8150 1.4050 ;
      RECT 3.9700 0.4250 4.1400 0.4800 ;
      RECT 7.2650 1.6450 7.9200 1.7350 ;
      RECT 7.8300 1.3650 7.9200 1.6450 ;
      RECT 7.4700 0.6100 7.9200 0.7000 ;
      RECT 7.8300 0.4450 7.9200 0.6100 ;
      RECT 7.4700 0.7000 7.5600 1.6450 ;
      RECT 3.9850 1.8300 7.3550 1.9200 ;
      RECT 7.2650 1.7350 7.3550 1.8300 ;
      RECT 4.9000 1.4950 4.9900 1.8300 ;
      RECT 4.9000 1.3250 5.0400 1.4950 ;
      RECT 0.5900 1.3200 0.7300 1.5150 ;
      RECT 0.6400 0.6900 0.7300 1.3200 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0450 1.6850 0.9100 1.7750 ;
      RECT 0.8200 1.0350 0.9100 1.6850 ;
      RECT 0.2550 0.8750 0.3450 1.6850 ;
      RECT 0.0950 0.7850 0.3450 0.8750 ;
      RECT 0.0950 0.4850 0.1850 0.7850 ;
      RECT 1.2600 0.7550 1.3500 1.8650 ;
      RECT 1.1550 0.6650 1.3500 0.7550 ;
      RECT 1.8050 1.4550 1.9450 1.8850 ;
      RECT 1.8550 0.6750 1.9450 1.4550 ;
      RECT 1.8100 0.5700 1.9450 0.6750 ;
      RECT 0.8900 0.4800 1.9450 0.5700 ;
      RECT 0.8900 0.5700 0.9800 0.8250 ;
      RECT 0.8900 0.8250 1.0900 0.9150 ;
      RECT 1.0000 0.9150 1.0900 1.8450 ;
      RECT 2.9100 1.7600 3.0000 1.9800 ;
      RECT 2.2500 1.6700 3.0000 1.7600 ;
      RECT 2.2500 0.8250 3.1650 0.9150 ;
      RECT 2.2500 0.9150 2.3400 1.6700 ;
  END
END M2SDFFQ_X3M_A12TH

MACRO M2SDFFQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6800 ;
        RECT 2.6150 0.3200 2.7850 0.5250 ;
        RECT 3.2350 0.3200 3.4050 0.5300 ;
        RECT 4.9150 0.3200 5.0850 0.3850 ;
        RECT 8.3300 0.3200 8.5000 0.4600 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7550 1.2500 3.2050 1.3500 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0500 2.8750 1.1500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.6400 0.8350 8.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.8150 7.5500 1.2500 ;
        RECT 7.0600 1.2500 7.6750 1.3500 ;
        RECT 7.0000 0.7150 7.7100 0.8150 ;
        RECT 7.0600 1.3500 7.1500 1.7200 ;
        RECT 7.5750 1.3500 7.6750 1.7250 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 4.3800 2.0500 4.5500 2.0800 ;
        RECT 0.3150 1.8750 0.4850 2.0800 ;
        RECT 8.3100 1.8400 8.4800 2.0800 ;
        RECT 2.6650 1.8000 2.7650 2.0800 ;
        RECT 3.2550 1.6350 3.3650 2.0800 ;
        RECT 1.5350 1.5700 1.6350 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 0.5900 1.3200 0.7300 1.5150 ;
      RECT 0.6400 0.5550 0.7300 1.3200 ;
      RECT 0.0450 1.6750 0.9100 1.7650 ;
      RECT 0.8200 1.0350 0.9100 1.6750 ;
      RECT 0.2550 0.8750 0.3450 1.6750 ;
      RECT 0.0950 0.7850 0.3450 0.8750 ;
      RECT 0.0950 0.5550 0.1850 0.7850 ;
      RECT 1.2600 0.7550 1.3500 1.8450 ;
      RECT 1.1750 0.6650 1.3500 0.7550 ;
      RECT 0.9000 0.4800 1.9000 0.5700 ;
      RECT 1.8100 0.5700 1.9000 1.8850 ;
      RECT 1.0000 0.9150 1.0900 1.8450 ;
      RECT 0.9000 0.8250 1.0900 0.9150 ;
      RECT 0.9000 0.5700 0.9900 0.8250 ;
      RECT 2.2500 1.5250 3.1500 1.6150 ;
      RECT 2.2500 0.8250 3.1650 0.9150 ;
      RECT 2.2500 0.9150 2.3400 1.5250 ;
      RECT 2.0700 0.6250 3.4250 0.7150 ;
      RECT 3.3350 0.7150 3.4250 1.2950 ;
      RECT 2.0700 0.7150 2.1600 1.8850 ;
      RECT 2.0700 0.5000 2.1600 0.6250 ;
      RECT 3.5350 0.4650 3.6250 1.9000 ;
      RECT 3.8000 1.6200 3.8900 1.9400 ;
      RECT 3.8000 1.5300 4.0100 1.6200 ;
      RECT 3.9200 1.1300 4.0100 1.5300 ;
      RECT 3.9200 1.0400 5.0550 1.1300 ;
      RECT 3.9200 0.6800 4.0100 1.0400 ;
      RECT 4.2900 1.6000 5.3200 1.6900 ;
      RECT 4.2900 1.2550 4.3800 1.6000 ;
      RECT 5.2300 0.7750 5.3200 1.6000 ;
      RECT 4.6550 0.6850 5.3200 0.7750 ;
      RECT 6.1800 1.5750 6.7050 1.6650 ;
      RECT 6.1800 1.3050 6.2700 1.5750 ;
      RECT 6.6150 0.9550 6.7050 1.5750 ;
      RECT 6.5150 0.8650 6.7050 0.9550 ;
      RECT 6.8000 1.0700 7.3400 1.1600 ;
      RECT 5.6150 1.6400 5.7050 1.7200 ;
      RECT 5.6150 1.5500 6.0900 1.6400 ;
      RECT 6.0000 1.1900 6.0900 1.5500 ;
      RECT 6.0000 1.1000 6.5000 1.1900 ;
      RECT 6.0000 0.7700 6.0900 1.1000 ;
      RECT 5.6100 0.6800 6.8900 0.7700 ;
      RECT 5.6100 0.7700 5.7000 0.8350 ;
      RECT 6.8000 0.7700 6.8900 1.0700 ;
      RECT 5.6100 0.6650 5.7000 0.6800 ;
      RECT 3.7400 0.4800 8.1800 0.5700 ;
      RECT 8.0900 0.5700 8.1800 1.5300 ;
      RECT 5.8200 1.1650 5.9100 1.4400 ;
      RECT 5.4100 1.0750 5.9100 1.1650 ;
      RECT 5.4100 0.5700 5.5000 1.0750 ;
      RECT 3.7400 0.5700 3.8300 1.4200 ;
      RECT 3.9850 0.4250 4.1550 0.4800 ;
      RECT 8.0750 1.6450 8.7200 1.7350 ;
      RECT 8.6300 1.3650 8.7200 1.6450 ;
      RECT 8.2750 0.6100 8.7200 0.7000 ;
      RECT 8.6300 0.4450 8.7200 0.6100 ;
      RECT 8.2750 0.7000 8.3650 1.6450 ;
      RECT 4.0400 1.8300 8.1650 1.9200 ;
      RECT 8.0750 1.7350 8.1650 1.8300 ;
      RECT 4.0400 1.7300 4.1300 1.8300 ;
      RECT 5.4350 1.3900 5.5250 1.8300 ;
      RECT 5.4350 1.3000 5.6250 1.3900 ;
  END
END M2SDFFQ_X4M_A12TH

MACRO MX2_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.6250 0.3200 0.7400 0.6800 ;
        RECT 1.9150 0.3200 2.0850 0.7000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7900 1.1500 1.3000 ;
        RECT 0.8950 1.3000 1.1500 1.4000 ;
        RECT 1.0500 0.6900 1.3100 0.7900 ;
        RECT 0.8950 1.4000 0.9950 1.7300 ;
    END
    ANTENNADIFFAREA 0.151 ;
  END Y

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.5800 0.9500 1.0000 ;
        RECT 0.5450 1.0000 0.9500 1.1000 ;
        RECT 0.8500 0.4800 1.7150 0.5800 ;
        RECT 0.5450 0.9100 0.6350 1.0000 ;
        RECT 1.6150 0.5800 1.7150 0.8000 ;
        RECT 1.6150 0.8000 2.1200 0.9000 ;
        RECT 2.0300 0.9000 2.1200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0650 1.7650 0.1850 2.0800 ;
        RECT 0.6350 1.7600 0.7350 2.0800 ;
        RECT 1.1550 1.7600 1.2550 2.0800 ;
        RECT 1.4150 1.7300 1.5050 2.0800 ;
        RECT 1.9550 1.7100 2.0650 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1900 0.1500 1.4850 ;
        RECT 0.0500 1.0900 0.2350 1.1900 ;
    END
    ANTENNAGATEAREA 0.0273 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 1.0100 1.7500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0273 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.3350 1.3300 0.7950 1.4200 ;
      RECT 0.7050 1.2100 0.7950 1.3300 ;
      RECT 0.3350 1.4200 0.4350 1.9750 ;
      RECT 0.3350 0.8600 0.4250 1.3300 ;
      RECT 0.0800 0.7700 0.4250 0.8600 ;
      RECT 0.0800 0.6500 0.1700 0.7700 ;
      RECT 1.6700 1.6300 1.7700 1.9200 ;
      RECT 1.4150 1.5400 1.7700 1.6300 ;
      RECT 1.4150 1.1600 1.5050 1.5400 ;
      RECT 1.2400 1.0700 1.5050 1.1600 ;
      RECT 1.4150 0.6950 1.5050 1.0700 ;
      RECT 2.2300 1.5300 2.3200 1.7650 ;
      RECT 1.8900 1.4400 2.3200 1.5300 ;
      RECT 2.2300 0.6800 2.3200 1.4400 ;
      RECT 1.8900 1.3000 1.9800 1.4400 ;
  END
END MX2_X0P5B_A12TH

MACRO MX2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3450 0.3200 0.4450 0.7600 ;
        RECT 1.5100 0.3200 1.6800 0.5500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0700 0.8500 1.3900 0.9500 ;
        RECT 1.0700 0.9500 1.2950 0.9550 ;
        RECT 1.0700 0.6800 1.1650 0.8500 ;
        RECT 1.1950 0.9550 1.2950 1.9900 ;
    END
    ANTENNADIFFAREA 0.129375 ;
  END Y

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9500 0.3500 1.1900 ;
        RECT 0.2400 0.8500 0.6550 0.9500 ;
        RECT 0.5550 0.5700 0.6550 0.8500 ;
        RECT 0.5550 0.4800 1.3900 0.5700 ;
        RECT 1.3000 0.5700 1.3900 0.6500 ;
        RECT 1.3000 0.6500 1.7550 0.7400 ;
        RECT 1.6500 0.7400 1.7550 1.1100 ;
    END
    ANTENNAGATEAREA 0.0558 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.1850 0.7900 1.5700 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1650 1.9500 1.5900 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.4150 1.9350 1.5850 2.0800 ;
        RECT 0.9300 1.8600 1.0300 2.0800 ;
        RECT 2.0250 1.8600 2.1250 2.0800 ;
        RECT 0.3400 1.7200 0.4400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0600 1.2800 0.5300 1.3700 ;
      RECT 0.4400 1.3700 0.5300 1.4800 ;
      RECT 0.0600 1.7650 0.1950 1.9650 ;
      RECT 0.0600 1.3700 0.1500 1.7650 ;
      RECT 0.0600 0.7750 0.1500 1.2800 ;
      RECT 0.0600 0.6050 0.1900 0.7750 ;
      RECT 0.6100 1.7700 0.7100 1.8900 ;
      RECT 0.6100 1.6800 0.9800 1.7700 ;
      RECT 0.7650 0.6750 0.9800 0.7700 ;
      RECT 0.8900 1.2800 0.9800 1.6800 ;
      RECT 0.8900 0.7700 0.9800 1.0700 ;
      RECT 0.8900 1.0700 1.1050 1.2800 ;
      RECT 1.4100 1.6800 2.1500 1.7700 ;
      RECT 2.0600 0.6200 2.1500 1.6800 ;
      RECT 2.0100 0.4500 2.1500 0.6200 ;
      RECT 1.7650 1.7700 1.8650 1.9900 ;
      RECT 1.4100 1.4800 1.5000 1.6800 ;
  END
END MX2_X0P5M_A12TH

MACRO MX2_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.6250 0.3200 0.7400 0.5150 ;
        RECT 1.9450 0.3200 2.0650 0.6100 ;
    END
  END VSS

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5400 0.6500 0.9500 0.7500 ;
        RECT 0.8500 0.5800 0.9500 0.6500 ;
        RECT 0.5400 0.7500 0.6400 1.1350 ;
        RECT 0.8500 0.4800 1.7500 0.5800 ;
        RECT 1.6500 0.5800 1.7500 0.7000 ;
        RECT 1.6500 0.7000 2.1200 0.7900 ;
        RECT 2.0300 0.7900 2.1200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.6400 1.7300 0.7300 2.0800 ;
        RECT 1.1600 1.7300 1.2500 2.0800 ;
        RECT 1.4300 1.7050 1.5200 2.0800 ;
        RECT 1.9550 1.7050 2.0650 2.0800 ;
        RECT 0.0800 1.5950 0.1700 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1900 0.1500 1.4200 ;
        RECT 0.0500 1.0900 0.2400 1.1900 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7900 1.1500 1.2500 ;
        RECT 0.8950 1.2500 1.1500 1.3500 ;
        RECT 1.0500 0.6900 1.3100 0.7900 ;
        RECT 0.8950 1.3500 0.9950 1.9500 ;
    END
    ANTENNADIFFAREA 0.218875 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 1.0100 1.7500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.3400 1.3550 0.7950 1.4450 ;
      RECT 0.7050 1.2350 0.7950 1.3550 ;
      RECT 0.3400 1.4450 0.4300 1.7550 ;
      RECT 0.3400 0.9000 0.4300 1.3550 ;
      RECT 0.0800 0.8100 0.4300 0.9000 ;
      RECT 0.0800 0.6350 0.1700 0.8100 ;
      RECT 1.6850 1.5900 1.7850 1.8750 ;
      RECT 1.4300 1.5000 1.7850 1.5900 ;
      RECT 1.4300 1.1600 1.5200 1.5000 ;
      RECT 1.2400 1.0700 1.5200 1.1600 ;
      RECT 1.4300 0.6800 1.5200 1.0700 ;
      RECT 2.2300 1.4700 2.3200 1.9400 ;
      RECT 1.8900 1.3800 2.3200 1.4700 ;
      RECT 2.2300 0.6800 2.3200 1.3800 ;
      RECT 1.8900 1.2400 1.9800 1.3800 ;
  END
END MX2_X0P7B_A12TH

MACRO MX2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7400 ;
        RECT 1.5050 0.3200 1.6750 0.4250 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0700 0.8500 1.3900 0.9500 ;
        RECT 1.0700 0.9500 1.2950 0.9550 ;
        RECT 1.0700 0.7150 1.1700 0.8500 ;
        RECT 1.1950 0.9550 1.2950 1.9900 ;
    END
    ANTENNADIFFAREA 0.1805 ;
  END Y

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9500 0.3500 1.1900 ;
        RECT 0.2400 0.8500 0.6550 0.9500 ;
        RECT 0.5550 0.6050 0.6550 0.8500 ;
        RECT 0.5550 0.5150 1.7550 0.6050 ;
        RECT 1.6500 0.6050 1.7550 1.1100 ;
    END
    ANTENNAGATEAREA 0.0777 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0600 0.7900 1.5000 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1650 1.9500 1.5900 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.4150 1.9350 1.5850 2.0800 ;
        RECT 0.9300 1.8600 1.0300 2.0800 ;
        RECT 2.0250 1.8600 2.1250 2.0800 ;
        RECT 0.3400 1.5950 0.4400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0600 1.2800 0.5300 1.3700 ;
      RECT 0.4400 1.3700 0.5300 1.4800 ;
      RECT 0.0600 1.6000 0.2150 1.9800 ;
      RECT 0.0600 1.3700 0.1500 1.6000 ;
      RECT 0.0600 0.7600 0.1500 1.2800 ;
      RECT 0.0600 0.5500 0.1900 0.7600 ;
      RECT 0.5550 1.6800 0.9800 1.7700 ;
      RECT 0.7650 0.7250 0.9800 0.8200 ;
      RECT 0.8900 1.2800 0.9800 1.6800 ;
      RECT 0.8900 0.8200 0.9800 1.0700 ;
      RECT 0.8900 1.0700 1.1050 1.2800 ;
      RECT 1.4100 1.6800 2.1500 1.7700 ;
      RECT 2.0600 0.6800 2.1500 1.6800 ;
      RECT 2.0100 0.5100 2.1500 0.6800 ;
      RECT 1.7650 1.7700 1.8650 1.9500 ;
      RECT 1.4100 1.2800 1.5000 1.6800 ;
  END
END MX2_X0P7M_A12TH

MACRO MX2_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.6700 0.3200 0.7700 0.6300 ;
        RECT 2.0700 0.3200 2.1600 0.9400 ;
    END
  END VSS

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.5800 1.9500 1.0500 ;
        RECT 1.8500 1.0500 2.2750 1.1600 ;
        RECT 0.8600 0.4800 1.9500 0.5800 ;
        RECT 0.8600 0.5800 0.9600 0.8000 ;
        RECT 0.5550 0.8000 0.9600 0.9000 ;
        RECT 0.5550 0.9000 0.6450 1.2350 ;
    END
    ANTENNAGATEAREA 0.0954 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.7050 1.7900 0.7950 2.0800 ;
        RECT 1.5000 1.7900 1.6200 2.0800 ;
        RECT 1.2250 1.7700 1.3150 2.0800 ;
        RECT 2.1000 1.5700 2.1900 2.0800 ;
        RECT 0.0950 1.5000 0.2150 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1500 0.1500 1.3900 ;
        RECT 0.0500 1.0400 0.2350 1.1500 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9200 1.1500 1.3050 ;
        RECT 0.9650 1.3050 1.1500 1.4050 ;
        RECT 1.0500 0.8050 1.3600 0.9200 ;
        RECT 0.9650 1.4050 1.0550 1.7500 ;
    END
    ANTENNADIFFAREA 0.317 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.0100 1.7600 1.4550 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.3700 1.3600 0.8750 1.4500 ;
      RECT 0.7850 1.0250 0.8750 1.3600 ;
      RECT 0.3700 1.4500 0.4600 1.6900 ;
      RECT 0.3700 0.8900 0.4600 1.3600 ;
      RECT 0.0500 0.8000 0.4600 0.8900 ;
      RECT 1.7700 1.6850 1.8700 1.9850 ;
      RECT 1.4550 1.5950 1.8700 1.6850 ;
      RECT 1.4550 0.7900 1.6650 0.9000 ;
      RECT 1.4550 1.1850 1.5450 1.5950 ;
      RECT 1.2700 1.0600 1.5450 1.1850 ;
      RECT 1.4550 0.9000 1.5450 1.0600 ;
      RECT 2.3650 1.4200 2.4550 1.9600 ;
      RECT 1.9300 1.3300 2.4550 1.4200 ;
      RECT 2.3650 0.7500 2.4550 1.3300 ;
  END
END MX2_X1B_A12TH

MACRO MX2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7400 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1950 1.9500 1.6300 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0700 0.8500 1.3900 0.9500 ;
        RECT 1.0700 0.9500 1.2950 0.9550 ;
        RECT 1.0700 0.7050 1.1700 0.8500 ;
        RECT 1.1950 0.9550 1.2950 1.9900 ;
    END
    ANTENNADIFFAREA 0.2472 ;
  END Y

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9500 0.3500 1.1900 ;
        RECT 0.2400 0.8500 0.6550 0.9500 ;
        RECT 0.5550 0.5800 0.6550 0.8500 ;
        RECT 0.5550 0.4800 1.7600 0.5800 ;
        RECT 1.6600 0.5800 1.7600 1.2800 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0600 0.7900 1.5900 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.4500 1.9400 1.5500 2.0800 ;
        RECT 2.0250 1.9200 2.1250 2.0800 ;
        RECT 0.9300 1.8800 1.0300 2.0800 ;
        RECT 0.3400 1.5600 0.4400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0600 1.2800 0.5300 1.3700 ;
      RECT 0.4400 1.3700 0.5300 1.4600 ;
      RECT 0.0600 1.5750 0.2150 1.9550 ;
      RECT 0.0600 1.3700 0.1500 1.5750 ;
      RECT 0.0600 0.7600 0.1500 1.2800 ;
      RECT 0.0600 0.5500 0.1900 0.7600 ;
      RECT 0.6150 1.7700 0.7100 1.8850 ;
      RECT 0.6150 1.6800 0.9800 1.7700 ;
      RECT 0.7450 0.7000 0.9800 0.7950 ;
      RECT 0.8900 1.2800 0.9800 1.6800 ;
      RECT 0.8900 0.7950 0.9800 1.0700 ;
      RECT 0.8900 1.0700 1.1050 1.2800 ;
      RECT 1.4100 1.7400 2.1450 1.8300 ;
      RECT 2.0550 0.9700 2.1450 1.7400 ;
      RECT 2.0050 0.7600 2.1450 0.9700 ;
      RECT 1.7650 1.8300 1.8650 1.9500 ;
      RECT 1.4100 1.2700 1.5000 1.7400 ;
  END
END MX2_X1M_A12TH

MACRO MX2_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.5750 0.3200 0.6750 0.7200 ;
        RECT 1.6100 0.3200 1.7800 0.3900 ;
        RECT 2.5650 0.3200 2.6650 0.5950 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9300 1.4500 2.7500 1.5500 ;
        RECT 1.9300 1.5500 2.0200 1.5900 ;
        RECT 2.3650 1.5500 2.4650 1.8800 ;
        RECT 2.6500 0.8050 2.7500 1.4500 ;
        RECT 1.8100 1.5900 2.0200 1.6800 ;
        RECT 2.0700 0.7050 2.7500 0.8050 ;
        RECT 1.8100 1.6800 1.9800 1.8800 ;
        RECT 2.0700 0.4550 2.2400 0.7050 ;
    END
    ANTENNADIFFAREA 0.365 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0300 0.8500 1.4150 0.9600 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0600 0.7600 1.2400 ;
        RECT 0.5550 0.8500 0.7600 1.0600 ;
    END
    ANTENNAGATEAREA 0.1197 ;
  END S0

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.8100 0.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.5050 2.0100 0.6750 2.0800 ;
        RECT 0.9850 2.0100 1.1550 2.0800 ;
        RECT 1.5400 2.0100 1.7100 2.0800 ;
        RECT 0.1100 1.9700 0.2100 2.0800 ;
        RECT 2.1100 1.6600 2.2050 2.0800 ;
        RECT 2.6250 1.6600 2.7250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8500 1.0500 1.4600 1.1400 ;
      RECT 0.8300 1.3000 0.9400 1.7200 ;
      RECT 0.8500 1.1400 0.9400 1.3000 ;
      RECT 0.8500 0.4100 0.9400 1.0500 ;
      RECT 1.5700 0.9250 2.3550 1.0150 ;
      RECT 1.2700 1.4500 1.4400 1.7400 ;
      RECT 1.3500 1.3200 1.4400 1.4500 ;
      RECT 1.3500 1.2300 1.6600 1.3200 ;
      RECT 1.5700 1.0150 1.6600 1.2300 ;
      RECT 1.5700 0.5700 1.6600 0.9250 ;
      RECT 1.1300 0.4800 1.6600 0.5700 ;
      RECT 1.7500 1.2450 2.5550 1.3350 ;
      RECT 2.4650 1.1250 2.5550 1.2450 ;
      RECT 0.3300 1.8300 1.6200 1.9200 ;
      RECT 1.5300 1.5000 1.6200 1.8300 ;
      RECT 1.5300 1.4100 1.8400 1.5000 ;
      RECT 1.7500 1.3350 1.8400 1.4100 ;
      RECT 1.7500 1.1250 1.8400 1.2450 ;
      RECT 0.3300 1.5300 0.4200 1.8300 ;
      RECT 0.0450 1.4400 0.4200 1.5300 ;
      RECT 0.0450 0.7000 0.1350 1.4400 ;
      RECT 0.0450 0.6100 0.2200 0.7000 ;
      RECT 0.1300 0.4900 0.2200 0.6100 ;
  END
END MX2_X1P4B_A12TH

MACRO MX2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7250 ;
        RECT 0.9550 0.3200 1.1250 0.4150 ;
        RECT 2.1250 0.3200 2.2250 0.7500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.7700 1.0600 ;
        RECT 0.6800 1.0600 0.7700 1.6550 ;
        RECT 0.4500 0.7050 0.7700 0.8100 ;
    END
    ANTENNADIFFAREA 0.3137 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9100 1.5500 1.3300 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9100 1.2050 2.2800 1.3050 ;
        RECT 2.0100 1.3050 2.2800 1.3500 ;
    END
    ANTENNAGATEAREA 0.105 ;
  END S0

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.2800 2.7500 1.4100 ;
        RECT 2.5500 1.0700 2.7500 1.2800 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.0650 1.8000 1.1650 2.0800 ;
        RECT 0.2900 1.7700 0.3900 2.0800 ;
        RECT 1.5950 1.7250 1.6950 2.0800 ;
        RECT 2.6250 1.6800 2.7250 2.0800 ;
        RECT 2.1050 1.5000 2.2050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0650 0.6850 1.6050 0.7850 ;
      RECT 0.4800 1.7450 0.9700 1.8350 ;
      RECT 0.8800 1.6900 0.9700 1.7450 ;
      RECT 0.4800 1.2400 0.5700 1.7450 ;
      RECT 0.2000 1.1500 0.5700 1.2400 ;
      RECT 0.8800 1.6000 1.4300 1.6900 ;
      RECT 1.3400 1.6900 1.4300 1.9900 ;
      RECT 1.0650 0.7850 1.1550 1.6000 ;
      RECT 1.8500 1.5100 1.9400 1.8300 ;
      RECT 1.2450 1.4200 1.9400 1.5100 ;
      RECT 1.7300 0.7150 1.8200 1.4200 ;
      RECT 1.2450 1.2800 1.3350 1.4200 ;
      RECT 1.9300 0.8600 2.6700 0.9500 ;
      RECT 2.5800 0.5600 2.6700 0.8600 ;
      RECT 2.3700 0.9500 2.4600 1.8500 ;
      RECT 0.8650 0.5950 0.9550 1.1200 ;
      RECT 0.2700 0.5950 0.3600 0.9050 ;
      RECT 0.0950 0.9050 0.3600 1.0000 ;
      RECT 1.9300 0.5950 2.0200 0.8600 ;
      RECT 0.2700 0.5050 2.0200 0.5950 ;
  END
END MX2_X1P4M_A12TH

MACRO MX2_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.5650 0.3200 0.6750 0.3900 ;
        RECT 1.6100 0.3200 1.7200 0.3900 ;
        RECT 2.5650 0.3200 2.6650 0.6300 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8950 0.3500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8250 0.7500 1.2800 ;
    END
    ANTENNAGATEAREA 0.1554 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1450 0.8500 1.3900 0.9500 ;
        RECT 1.1450 0.9500 1.2350 1.1700 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.6500 2.7500 1.7500 ;
        RECT 1.8500 1.7500 1.9400 1.9900 ;
        RECT 2.3700 1.7500 2.4600 1.9900 ;
        RECT 1.8500 1.5600 1.9400 1.6500 ;
        RECT 2.6500 0.8200 2.7500 1.6500 ;
        RECT 2.1100 0.7300 2.7500 0.8200 ;
        RECT 2.1100 0.4500 2.2000 0.7300 ;
    END
    ANTENNADIFFAREA 0.518 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.0650 1.8400 1.1650 2.0800 ;
        RECT 2.1050 1.8400 2.2050 2.0800 ;
        RECT 2.6250 1.8400 2.7250 2.0800 ;
        RECT 1.5850 1.7700 1.6850 2.0800 ;
        RECT 0.5950 1.6000 0.6950 2.0800 ;
        RECT 0.0750 1.5300 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8600 1.2800 1.5050 1.3700 ;
      RECT 1.4150 1.1300 1.5050 1.2800 ;
      RECT 0.8600 1.3700 0.9500 1.7400 ;
      RECT 0.8600 0.7000 0.9500 1.2800 ;
      RECT 1.9550 1.0900 2.3450 1.1800 ;
      RECT 1.3300 1.5500 1.4200 1.9800 ;
      RECT 1.3300 1.4600 1.6850 1.5500 ;
      RECT 1.5950 1.3900 1.6850 1.4600 ;
      RECT 1.5950 0.7600 1.6850 1.3000 ;
      RECT 1.0750 0.6600 1.6850 0.7600 ;
      RECT 1.5950 1.3000 2.0450 1.3900 ;
      RECT 1.9550 1.1800 2.0450 1.3000 ;
      RECT 1.7750 0.9100 2.5550 1.0000 ;
      RECT 2.4650 1.0000 2.5550 1.2100 ;
      RECT 0.4400 0.4800 1.8650 0.5700 ;
      RECT 1.7750 0.5700 1.8650 0.9100 ;
      RECT 1.7750 1.0000 1.8650 1.1900 ;
      RECT 0.3400 1.5000 0.4300 1.8400 ;
      RECT 0.3400 1.4100 0.5300 1.5000 ;
      RECT 0.4400 0.7800 0.5300 1.4100 ;
      RECT 0.1250 0.6900 0.5300 0.7800 ;
      RECT 0.4400 0.5700 0.5300 0.6900 ;
      RECT 0.1250 0.4100 0.2150 0.6900 ;
  END
END MX2_X2B_A12TH

MACRO MX2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.5600 0.3200 0.6550 0.7200 ;
        RECT 1.6550 0.3200 1.7550 0.4700 ;
        RECT 2.5750 0.3200 2.6750 0.6400 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2200 0.3500 1.3900 ;
        RECT 0.2100 1.0100 0.3500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0687 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0100 0.7500 1.5000 ;
    END
    ANTENNAGATEAREA 0.1356 ;
  END S0

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.5000 1.1500 1.7900 ;
        RECT 1.0500 1.3300 1.2250 1.5000 ;
    END
    ANTENNAGATEAREA 0.0687 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.6500 2.7550 1.7500 ;
        RECT 1.8500 1.7500 1.9400 1.9900 ;
        RECT 2.3700 1.7500 2.4600 1.9900 ;
        RECT 1.8500 1.5900 1.9400 1.6500 ;
        RECT 2.6550 0.9800 2.7550 1.6500 ;
        RECT 2.1200 0.8900 2.7550 0.9800 ;
        RECT 2.1200 0.5400 2.2100 0.8900 ;
    END
    ANTENNADIFFAREA 0.402 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.1050 1.8400 2.2050 2.0800 ;
        RECT 2.6250 1.8400 2.7250 2.0800 ;
        RECT 1.5850 1.8200 1.6850 2.0800 ;
        RECT 0.5950 1.6600 0.6950 2.0800 ;
        RECT 0.0750 1.5900 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8600 1.0850 1.4950 1.1850 ;
      RECT 1.4000 1.1850 1.4950 1.2950 ;
      RECT 0.8600 1.1850 0.9500 1.8200 ;
      RECT 0.9450 0.6900 1.0350 1.0850 ;
      RECT 1.5850 1.3500 2.3650 1.4400 ;
      RECT 1.3300 1.6900 1.4200 1.9900 ;
      RECT 1.1950 0.6600 1.2850 0.7700 ;
      RECT 1.3300 1.6000 1.6850 1.6900 ;
      RECT 1.5850 1.4400 1.6850 1.6000 ;
      RECT 1.5850 0.8600 1.6750 1.3500 ;
      RECT 1.1950 0.7700 1.6750 0.8600 ;
      RECT 1.7650 1.0700 2.5650 1.1600 ;
      RECT 2.4750 1.1600 2.5650 1.2800 ;
      RECT 0.7650 0.4800 1.5350 0.5600 ;
      RECT 0.1150 0.8100 0.8550 0.9000 ;
      RECT 0.7650 0.5700 0.8550 0.8100 ;
      RECT 0.7650 0.5600 1.8550 0.5700 ;
      RECT 1.4450 0.5700 1.8550 0.6500 ;
      RECT 1.7650 0.6500 1.8550 1.0700 ;
      RECT 1.7650 1.1600 1.8550 1.2400 ;
      RECT 0.3400 1.5700 0.4300 1.9150 ;
      RECT 0.3400 1.4800 0.5500 1.5700 ;
      RECT 0.4600 0.9000 0.5500 1.4800 ;
      RECT 0.1150 0.4700 0.2050 0.8100 ;
  END
END MX2_X2M_A12TH

MACRO MX2_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6700 ;
        RECT 1.0700 0.3200 1.2600 0.5550 ;
        RECT 1.5750 0.3200 1.7650 0.5550 ;
        RECT 2.6200 0.3200 2.8100 0.5550 ;
        RECT 3.7050 0.3200 3.8050 0.6250 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5400 1.0500 0.9850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1188 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9650 1.2500 2.5150 1.3500 ;
    END
    ANTENNAGATEAREA 0.1188 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 1.0500 2.6350 1.1500 ;
    END
    ANTENNAGATEAREA 0.2154 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 1.6250 1.7600 1.7250 2.0800 ;
        RECT 2.1450 1.7600 2.2450 2.0800 ;
        RECT 2.6650 1.7600 2.7650 2.0800 ;
        RECT 3.1850 1.7500 3.2850 2.0800 ;
        RECT 3.7050 1.7500 3.8050 2.0800 ;
        RECT 4.2250 1.7500 4.3250 2.0800 ;
        RECT 0.0750 1.7350 0.1750 2.0800 ;
        RECT 0.5950 1.7350 0.6950 2.0800 ;
        RECT 1.1150 1.7350 1.2150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9250 1.4500 4.3500 1.5500 ;
        RECT 2.9250 1.5500 3.0250 1.8900 ;
        RECT 3.4450 1.5500 3.5450 1.8900 ;
        RECT 3.9650 1.5500 4.0650 1.8900 ;
        RECT 4.2500 0.8400 4.3500 1.4500 ;
        RECT 3.1850 0.7500 4.3500 0.8400 ;
        RECT 3.1850 0.4300 3.2850 0.7500 ;
        RECT 4.2300 0.4300 4.3500 0.7500 ;
    END
    ANTENNADIFFAREA 0.816 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.3800 1.4000 1.4700 1.7400 ;
      RECT 0.2600 1.3000 1.4700 1.4000 ;
      RECT 1.3200 0.9400 1.4100 1.3000 ;
      RECT 1.3200 0.8500 1.5300 0.9400 ;
      RECT 0.2600 1.1550 0.3600 1.3000 ;
      RECT 2.7450 1.2100 3.9150 1.3000 ;
      RECT 3.5450 1.1200 3.9150 1.2100 ;
      RECT 1.8850 1.5900 1.9850 1.9400 ;
      RECT 2.4050 1.5900 2.5050 1.9400 ;
      RECT 1.8850 1.5000 2.8350 1.5900 ;
      RECT 2.7450 1.3000 2.8350 1.5000 ;
      RECT 2.7450 0.9350 2.8350 1.2100 ;
      RECT 2.0900 0.8450 2.8350 0.9350 ;
      RECT 2.9600 0.9400 4.1350 1.0300 ;
      RECT 4.0450 1.0300 4.1350 1.2350 ;
      RECT 0.3350 1.5900 0.4350 1.9400 ;
      RECT 0.0550 0.9350 0.1450 1.5000 ;
      RECT 0.0550 1.5000 0.9550 1.5900 ;
      RECT 0.8550 1.5900 0.9550 1.9400 ;
      RECT 0.0550 0.8450 0.7050 0.9350 ;
      RECT 0.5950 0.7550 0.7050 0.8450 ;
      RECT 0.5950 0.5050 0.6950 0.6650 ;
      RECT 0.5950 0.6650 3.0500 0.7550 ;
      RECT 2.9600 0.7550 3.0500 0.9400 ;
      RECT 2.9600 1.0300 3.3950 1.1200 ;
  END
END MX2_X3B_A12TH

MACRO MX2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.5200 ;
        RECT 1.1350 0.3200 1.2350 0.5500 ;
        RECT 2.4950 0.3200 2.5950 0.6250 ;
        RECT 3.5600 0.3200 3.6600 0.6250 ;
    END
  END VSS

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0150 1.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.1842 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.0900 1.7750 0.1900 2.0800 ;
        RECT 0.6100 1.7650 0.7100 2.0800 ;
        RECT 1.6700 1.7350 1.7700 2.0800 ;
        RECT 1.1350 1.6950 1.2350 2.0800 ;
        RECT 2.4950 1.6550 2.5950 2.0800 ;
        RECT 3.0400 1.6550 3.1400 2.0800 ;
        RECT 3.5600 1.6550 3.6600 2.0800 ;
        RECT 1.9500 1.6150 2.0500 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 1.4500 3.6750 1.5500 ;
        RECT 2.2100 1.5500 2.3100 1.9100 ;
        RECT 2.7800 1.5500 2.8800 1.9100 ;
        RECT 3.3000 1.5500 3.4000 1.9100 ;
        RECT 3.5750 0.8400 3.6750 1.4500 ;
        RECT 2.2200 0.7500 3.6750 0.8400 ;
        RECT 2.2200 0.5700 2.3100 0.7500 ;
        RECT 3.0400 0.4300 3.1400 0.7500 ;
        RECT 1.8950 0.4800 2.3100 0.5700 ;
    END
    ANTENNADIFFAREA 0.66075 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1000 0.6600 1.1900 ;
        RECT 0.4500 0.8400 0.5500 1.1000 ;
    END
    ANTENNAGATEAREA 0.0972 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0150 1.5850 1.4350 ;
    END
    ANTENNAGATEAREA 0.0972 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.8200 1.4900 0.9700 1.9100 ;
      RECT 0.8200 1.4600 0.9100 1.4900 ;
      RECT 0.2550 1.3600 0.9100 1.4600 ;
      RECT 0.8200 0.9300 0.9100 1.3600 ;
      RECT 0.8200 0.8400 1.0200 0.9300 ;
      RECT 0.2550 1.0450 0.3550 1.3600 ;
      RECT 1.9700 1.0550 3.2700 1.1450 ;
      RECT 0.3500 1.6400 0.4500 1.9900 ;
      RECT 0.0700 1.5500 0.4500 1.6400 ;
      RECT 0.0700 0.7500 0.1600 1.5500 ;
      RECT 0.5750 0.4150 0.7450 0.6600 ;
      RECT 0.0700 0.6600 2.0600 0.7500 ;
      RECT 1.9700 0.7500 2.0600 1.0550 ;
      RECT 1.7350 1.2550 3.4700 1.3450 ;
      RECT 3.3800 1.0250 3.4700 1.2550 ;
      RECT 1.4100 1.6150 1.5100 1.9750 ;
      RECT 1.4100 1.5250 1.8250 1.6150 ;
      RECT 1.7350 1.3450 1.8250 1.5250 ;
      RECT 1.7350 0.9300 1.8250 1.2550 ;
      RECT 1.6200 0.8400 1.8250 0.9300 ;
  END
END MX2_X3M_A12TH

MACRO MX2_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7350 ;
        RECT 1.1150 0.3200 1.2150 0.4850 ;
        RECT 1.6950 0.3200 1.7950 0.4850 ;
        RECT 2.7350 0.3200 2.8350 0.4850 ;
        RECT 3.7750 0.3200 3.8750 0.6400 ;
        RECT 4.8150 0.3200 4.9150 0.6500 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.0500 0.9850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1554 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0350 1.2500 2.5850 1.3500 ;
    END
    ANTENNAGATEAREA 0.1554 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5350 1.0500 2.7050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2766 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0750 1.7350 0.1750 2.0800 ;
        RECT 0.5950 1.7350 0.6950 2.0800 ;
        RECT 1.1150 1.7350 1.2150 2.0800 ;
        RECT 1.6950 1.7350 1.7950 2.0800 ;
        RECT 2.2150 1.7350 2.3150 2.0800 ;
        RECT 2.7350 1.7350 2.8350 2.0800 ;
        RECT 3.2550 1.7250 3.3550 2.0800 ;
        RECT 3.7750 1.7250 3.8750 2.0800 ;
        RECT 4.2950 1.7250 4.3950 2.0800 ;
        RECT 4.8150 1.7250 4.9150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9950 1.4500 4.9400 1.5500 ;
        RECT 2.9950 1.5500 3.0950 1.8800 ;
        RECT 3.5150 1.5500 3.6150 1.8800 ;
        RECT 4.0350 1.5500 4.1350 1.8800 ;
        RECT 4.5550 1.5500 4.6550 1.8800 ;
        RECT 4.8400 0.8400 4.9400 1.4500 ;
        RECT 3.2600 0.7500 4.9400 0.8400 ;
        RECT 3.2600 0.4300 3.3700 0.7500 ;
        RECT 4.2950 0.4300 4.3950 0.7500 ;
    END
    ANTENNADIFFAREA 0.948 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.3500 1.6150 1.5400 1.9050 ;
      RECT 1.3500 0.8500 1.5600 0.9400 ;
      RECT 1.3500 1.4000 1.4400 1.6150 ;
      RECT 0.2600 1.3000 1.4400 1.4000 ;
      RECT 1.3500 0.9400 1.4400 1.3000 ;
      RECT 0.2600 1.1550 0.3600 1.3000 ;
      RECT 4.1050 1.0450 4.5250 1.1400 ;
      RECT 3.3650 0.9300 4.2050 1.0200 ;
      RECT 4.1050 1.0200 4.2050 1.0450 ;
      RECT 0.3350 1.5900 0.4350 1.9900 ;
      RECT 0.0550 0.9350 0.1450 1.5000 ;
      RECT 0.0550 1.5000 0.9550 1.5900 ;
      RECT 0.8550 1.5900 0.9550 1.9900 ;
      RECT 0.0550 0.8450 0.7050 0.9350 ;
      RECT 0.5950 0.7550 0.7050 0.8450 ;
      RECT 0.5950 0.5050 0.6950 0.6650 ;
      RECT 0.5950 0.6650 3.1400 0.7550 ;
      RECT 3.0500 0.7550 3.1400 1.0500 ;
      RECT 3.0500 1.0500 3.4650 1.1400 ;
      RECT 3.3650 1.0200 3.4650 1.0500 ;
      RECT 3.8850 1.2300 4.7250 1.3200 ;
      RECT 4.6350 1.0250 4.7250 1.2300 ;
      RECT 1.9550 1.5900 2.0550 1.9900 ;
      RECT 2.4750 1.5900 2.5750 1.9900 ;
      RECT 1.9550 1.5000 2.9050 1.5900 ;
      RECT 2.8150 1.3200 2.9050 1.5000 ;
      RECT 2.8150 0.9350 2.9050 1.2300 ;
      RECT 2.1600 0.8450 2.9050 0.9350 ;
      RECT 2.8150 1.2300 3.6850 1.3200 ;
      RECT 3.5850 1.2100 3.6850 1.2300 ;
      RECT 3.5850 1.1200 3.9850 1.2100 ;
      RECT 3.8850 1.2100 3.9850 1.2300 ;
  END
END MX2_X4B_A12TH

MACRO MX2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6000 ;
        RECT 0.9950 0.3200 1.0950 0.6000 ;
        RECT 1.9100 0.3200 2.0800 0.5500 ;
        RECT 2.9300 0.3200 3.1000 0.5650 ;
        RECT 3.6700 0.3200 3.7700 0.8850 ;
        RECT 4.6250 0.3200 4.7250 0.8850 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3650 1.0400 2.8250 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9450 1.2500 4.3650 1.3500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1750 1.2500 3.1900 1.3500 ;
        RECT 2.1750 1.3500 2.2750 1.4700 ;
    END
    ANTENNAGATEAREA 0.2352 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6500 1.8400 1.7500 ;
        RECT 0.7100 1.7500 0.8000 1.9900 ;
        RECT 1.2300 1.7500 1.3200 1.9900 ;
        RECT 1.7500 1.7500 1.8400 1.9900 ;
        RECT 1.7500 1.5700 1.8400 1.6500 ;
        RECT 0.0500 0.7900 0.1500 1.6500 ;
        RECT 0.0500 0.6900 1.5850 0.7900 ;
        RECT 0.5350 0.4200 0.6350 0.6900 ;
        RECT 1.4850 0.4200 1.5850 0.6900 ;
    END
    ANTENNADIFFAREA 0.806 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.4450 1.8400 0.5450 2.0800 ;
        RECT 0.9650 1.8400 1.0650 2.0800 ;
        RECT 1.4850 1.8400 1.5850 2.0800 ;
        RECT 2.0050 1.8000 2.1050 2.0800 ;
        RECT 2.5250 1.8000 2.6250 2.0800 ;
        RECT 4.1050 1.8000 4.2050 2.0800 ;
        RECT 4.6250 1.8000 4.7250 2.0800 ;
        RECT 3.5750 1.7550 3.6750 2.0800 ;
        RECT 3.0450 1.7150 3.1450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.9950 1.5850 2.8800 1.6750 ;
      RECT 2.7900 1.6750 2.8800 1.9550 ;
      RECT 2.1650 0.8400 2.6350 0.9300 ;
      RECT 0.2450 1.2600 0.3350 1.3800 ;
      RECT 1.1300 1.2300 1.2300 1.3700 ;
      RECT 0.8400 1.1400 1.2300 1.2300 ;
      RECT 1.8550 1.1500 1.9550 1.3700 ;
      RECT 2.2700 1.6750 2.3600 1.9550 ;
      RECT 1.8550 1.0600 2.2550 1.1500 ;
      RECT 2.1650 0.9300 2.2550 1.0600 ;
      RECT 1.9950 1.4700 2.0850 1.5850 ;
      RECT 0.2450 1.3800 2.0850 1.4700 ;
      RECT 1.1300 1.3700 2.0850 1.3800 ;
      RECT 3.2950 1.4400 4.5650 1.5300 ;
      RECT 4.4750 1.3000 4.5650 1.4400 ;
      RECT 3.7450 1.3000 3.8350 1.4400 ;
      RECT 3.2950 1.5300 3.4000 1.9550 ;
      RECT 3.2950 0.9600 3.3850 1.4400 ;
      RECT 3.1950 0.8600 3.3850 0.9600 ;
      RECT 3.8500 1.6200 4.7450 1.7100 ;
      RECT 4.6550 1.0900 4.7450 1.6200 ;
      RECT 3.4750 1.0000 4.7450 1.0900 ;
      RECT 0.5100 0.9700 0.6150 1.2150 ;
      RECT 1.6150 0.9700 1.7150 1.1100 ;
      RECT 1.3250 1.1100 1.7150 1.2000 ;
      RECT 1.9500 0.7500 2.0400 0.8800 ;
      RECT 0.5100 0.8800 2.0400 0.9700 ;
      RECT 3.4750 0.7500 3.5650 1.0000 ;
      RECT 1.9500 0.6600 3.5650 0.7500 ;
      RECT 3.8500 1.7100 3.9400 1.9900 ;
      RECT 4.3700 1.7100 4.4600 1.9900 ;
      RECT 4.1250 0.6100 4.2150 1.0000 ;
  END
END MX2_X4M_A12TH

MACRO MX2_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.5850 0.3200 0.6850 0.5800 ;
        RECT 1.6200 0.3200 1.7200 0.5800 ;
        RECT 2.6050 0.3200 2.6950 0.6300 ;
        RECT 3.6450 0.3200 3.7350 0.6300 ;
        RECT 4.6700 0.3200 4.7600 0.6300 ;
        RECT 5.4800 0.3200 5.5700 0.4300 ;
        RECT 6.3750 0.3200 6.4750 0.6000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 0.8500 1.2850 0.9500 ;
        RECT 0.2300 0.9500 0.3300 1.2000 ;
        RECT 0.8950 0.9500 1.2850 1.0500 ;
    END
    ANTENNAGATEAREA 0.2286 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7950 1.0500 6.1450 1.1500 ;
        RECT 6.0550 1.0000 6.1450 1.0500 ;
        RECT 6.0550 0.9000 6.7700 1.0000 ;
        RECT 6.6700 1.0000 6.7700 1.4800 ;
    END
    ANTENNAGATEAREA 0.2286 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 1.0500 5.6850 1.1500 ;
        RECT 5.5850 1.1500 5.6850 1.2500 ;
        RECT 5.5850 1.2500 6.4100 1.3500 ;
        RECT 6.3100 1.1900 6.4100 1.2500 ;
        RECT 6.3100 1.0900 6.5200 1.1900 ;
    END
    ANTENNAGATEAREA 0.3978 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7650 1.4500 4.7700 1.5500 ;
        RECT 4.6800 0.8200 4.7700 1.4500 ;
        RECT 2.0850 0.7300 4.7700 0.8200 ;
        RECT 2.0850 0.4300 2.1850 0.7300 ;
        RECT 3.1250 0.4300 3.2150 0.7300 ;
        RECT 4.1650 0.4300 4.2550 0.7300 ;
    END
    ANTENNADIFFAREA 1.446 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 1.5600 1.8400 1.6600 2.0800 ;
        RECT 2.0800 1.8400 2.1800 2.0800 ;
        RECT 2.6000 1.8400 2.7000 2.0800 ;
        RECT 3.1200 1.8400 3.2200 2.0800 ;
        RECT 3.6400 1.8400 3.7400 2.0800 ;
        RECT 4.1600 1.8400 4.2600 2.0800 ;
        RECT 4.7750 1.8400 4.8750 2.0800 ;
        RECT 5.9250 1.7800 6.0250 2.0800 ;
        RECT 6.4450 1.7800 6.5450 2.0800 ;
        RECT 0.3300 1.7700 0.4200 2.0800 ;
        RECT 1.0300 1.7700 1.1200 2.0800 ;
        RECT 5.4050 1.7400 5.5050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0450 0.5500 0.1700 0.6700 ;
      RECT 0.0450 1.3400 1.3800 1.4300 ;
      RECT 0.0450 0.7600 0.1350 1.3400 ;
      RECT 0.0450 0.6700 1.9950 0.7600 ;
      RECT 0.6750 1.4300 0.7650 1.7700 ;
      RECT 1.0400 0.4400 1.2100 0.6700 ;
      RECT 1.2900 1.4300 1.3800 1.7700 ;
      RECT 1.9050 0.9100 4.1100 1.0000 ;
      RECT 1.9050 0.7600 1.9950 0.9100 ;
      RECT 4.0200 1.0400 4.3900 1.1300 ;
      RECT 4.0200 1.0000 4.1100 1.0400 ;
      RECT 1.9500 0.9100 2.3200 1.1300 ;
      RECT 2.9900 0.9100 3.3600 1.1300 ;
      RECT 1.7250 1.0300 1.8150 1.2200 ;
      RECT 1.7250 1.2200 4.5900 1.3100 ;
      RECT 4.5000 1.0300 4.5900 1.2200 ;
      RECT 2.4600 1.0900 2.8300 1.3100 ;
      RECT 3.5000 1.0900 3.8700 1.3100 ;
      RECT 5.0950 0.7050 5.3450 0.7950 ;
      RECT 1.4700 1.6600 5.2250 1.7500 ;
      RECT 5.0950 1.3400 5.2250 1.6600 ;
      RECT 5.0950 0.7950 5.1850 1.3400 ;
      RECT 1.4700 1.2300 1.5600 1.6600 ;
      RECT 0.5300 1.1400 1.5600 1.2300 ;
      RECT 1.4400 1.0100 1.5600 1.1400 ;
      RECT 5.6700 1.5900 6.9550 1.6800 ;
      RECT 6.8650 0.8000 6.9550 1.5900 ;
      RECT 5.9300 0.7100 6.9550 0.8000 ;
      RECT 6.8300 0.4100 6.9550 0.7100 ;
      RECT 4.8950 0.6150 4.9850 0.9200 ;
      RECT 4.8600 0.9200 4.9850 1.1300 ;
      RECT 5.6700 1.6800 5.7600 1.9600 ;
      RECT 5.9300 0.6150 6.0200 0.7100 ;
      RECT 4.8950 0.5250 6.0200 0.6150 ;
      RECT 5.9300 0.4100 6.0200 0.5250 ;
      RECT 6.1900 1.6800 6.2800 1.9600 ;
  END
END MX2_X6B_A12TH

MACRO MX2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6300 ;
        RECT 1.0050 0.3200 1.1050 0.6300 ;
        RECT 1.9450 0.3200 2.0450 0.6300 ;
        RECT 2.9250 0.3200 3.0250 0.5700 ;
        RECT 4.0250 0.3200 4.1250 0.5550 ;
        RECT 4.5950 0.3200 4.6950 0.5550 ;
        RECT 5.6300 0.3200 5.7200 0.6400 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3500 1.0500 3.7200 1.1900 ;
    END
    ANTENNAGATEAREA 0.1914 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9650 1.0500 5.3350 1.2000 ;
    END
    ANTENNAGATEAREA 0.1914 ;
  END A

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 1.0500 4.4150 1.1750 ;
        RECT 3.8500 1.1750 3.9500 1.3000 ;
        RECT 3.1450 1.3000 3.9500 1.3900 ;
        RECT 3.1450 1.0700 3.2350 1.3000 ;
    END
    ANTENNAGATEAREA 0.3414 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2050 1.6500 2.8250 1.7500 ;
        RECT 2.2050 1.7500 2.3050 1.9250 ;
        RECT 2.7250 1.7500 2.8250 1.9250 ;
        RECT 2.2050 1.5950 2.3050 1.6500 ;
        RECT 2.7250 1.5000 2.8250 1.6500 ;
        RECT 0.0650 1.4950 2.3050 1.5950 ;
        RECT 0.6450 1.5950 0.7450 1.9250 ;
        RECT 1.1650 1.5950 1.2650 1.9250 ;
        RECT 1.6850 1.5950 1.7850 1.9250 ;
        RECT 0.0650 0.8750 0.1650 1.4950 ;
        RECT 0.0650 0.7750 2.5650 0.8750 ;
        RECT 0.5350 0.4450 0.6350 0.7750 ;
        RECT 1.4850 0.4450 1.5850 0.7750 ;
        RECT 2.4600 0.4450 2.5650 0.7750 ;
    END
    ANTENNADIFFAREA 1.207 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 2.4650 1.8400 2.5650 2.0800 ;
        RECT 0.3850 1.7700 0.4850 2.0800 ;
        RECT 0.9050 1.7700 1.0050 2.0800 ;
        RECT 1.4250 1.7700 1.5250 2.0800 ;
        RECT 1.9450 1.7700 2.0450 2.0800 ;
        RECT 2.9850 1.7700 3.0850 2.0800 ;
        RECT 3.5050 1.7700 3.6050 2.0800 ;
        RECT 5.1050 1.7700 5.2050 2.0800 ;
        RECT 5.6250 1.7700 5.7250 2.0800 ;
        RECT 4.0400 1.6350 4.1400 2.0800 ;
        RECT 4.5800 1.6350 4.6800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.9650 1.5400 3.8600 1.6300 ;
      RECT 3.7700 1.6300 3.8600 1.9700 ;
      RECT 2.9650 0.8600 3.6400 0.9500 ;
      RECT 3.4700 0.6600 3.6400 0.8600 ;
      RECT 0.2650 1.1950 0.3550 1.2950 ;
      RECT 1.8050 1.2250 2.1750 1.2950 ;
      RECT 2.9650 1.3850 3.0550 1.5400 ;
      RECT 0.2650 1.2950 3.0550 1.3850 ;
      RECT 2.8350 1.1950 3.0550 1.2950 ;
      RECT 2.9650 0.9500 3.0550 1.1950 ;
      RECT 3.2500 1.6350 3.3400 1.9700 ;
      RECT 2.9650 1.6300 3.3400 1.6350 ;
      RECT 4.3150 1.3650 5.5650 1.4550 ;
      RECT 5.4750 1.0700 5.5650 1.3650 ;
      RECT 4.3150 1.4550 4.4050 1.7950 ;
      RECT 4.7450 0.9150 4.8350 1.3650 ;
      RECT 4.2550 0.8250 4.8350 0.9150 ;
      RECT 0.5950 0.9650 2.8750 1.0550 ;
      RECT 0.5950 1.0550 0.6850 1.2050 ;
      RECT 2.7850 0.7500 2.8750 0.9650 ;
      RECT 2.7850 0.6600 3.3800 0.7500 ;
      RECT 3.2900 0.5700 3.3800 0.6600 ;
      RECT 3.2900 0.4800 3.8200 0.5700 ;
      RECT 3.7300 0.5700 3.8200 0.6450 ;
      RECT 3.7300 0.6450 5.2000 0.7350 ;
      RECT 4.8500 1.6550 4.9400 1.9750 ;
      RECT 4.8500 1.5650 5.7450 1.6550 ;
      RECT 5.1100 0.4300 5.2000 0.6450 ;
      RECT 5.1100 0.7350 5.2000 0.7700 ;
      RECT 5.1100 0.7700 5.7450 0.8600 ;
      RECT 5.3700 1.6550 5.4600 1.9750 ;
      RECT 5.6550 0.8600 5.7450 1.5650 ;
      RECT 1.4150 0.9650 1.6250 1.2000 ;
      RECT 2.3250 0.9650 2.6950 1.2000 ;
  END
END MX2_X6M_A12TH

MACRO MX2_X8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.5850 ;
        RECT 1.1150 0.3200 1.2150 0.5850 ;
        RECT 2.1550 0.3200 2.2550 0.5850 ;
        RECT 3.1950 0.3200 3.2950 0.5850 ;
        RECT 4.2150 0.3200 4.3050 0.6350 ;
        RECT 5.2000 0.3200 5.2900 0.6350 ;
        RECT 6.1250 0.3200 6.2150 0.6350 ;
        RECT 6.6450 0.3200 6.7350 0.4500 ;
        RECT 7.7050 0.3200 7.8050 0.4500 ;
        RECT 8.6250 0.3200 8.7250 0.6700 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.7000 5.9500 0.9400 ;
        RECT 4.6150 0.9400 5.9500 1.0500 ;
    END
    ANTENNAGATEAREA 0.3036 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 1.0400 7.3500 1.3800 ;
        RECT 7.2500 1.3800 8.2750 1.4800 ;
        RECT 8.1850 1.0000 8.2750 1.3800 ;
    END
    ANTENNAGATEAREA 0.3036 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.4400 3.5650 1.5600 ;
        RECT 3.4450 1.5600 3.5650 1.8000 ;
        RECT 0.3250 1.5600 0.4450 1.8800 ;
        RECT 0.8450 1.5600 0.9650 1.8800 ;
        RECT 1.3650 1.5600 1.4850 1.8800 ;
        RECT 1.8850 1.5600 2.0050 1.8800 ;
        RECT 2.4050 1.5600 2.5250 1.8800 ;
        RECT 2.9250 1.5600 3.0450 1.8800 ;
        RECT 0.0450 0.7950 0.1650 1.4400 ;
        RECT 3.4450 1.8000 4.1300 1.9200 ;
        RECT 0.0450 0.6750 3.8250 0.7950 ;
        RECT 0.5850 0.4100 0.7050 0.6750 ;
        RECT 1.6250 0.4100 1.7450 0.6750 ;
        RECT 2.6650 0.4100 2.7850 0.6750 ;
        RECT 3.7050 0.4100 3.8250 0.6750 ;
    END
    ANTENNADIFFAREA 1.928 ;
  END Y

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0600 1.0450 6.4900 1.1550 ;
        RECT 6.0600 1.1550 6.1600 1.1650 ;
        RECT 4.3900 1.1650 6.1600 1.2650 ;
        RECT 4.3900 1.0650 4.4950 1.1650 ;
    END
    ANTENNAGATEAREA 0.4968 ;
  END S0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 3.7200 2.0100 3.8100 2.0800 ;
        RECT 4.2350 1.8200 4.3350 2.0800 ;
        RECT 4.7550 1.8200 4.8550 2.0800 ;
        RECT 5.2750 1.8200 5.3750 2.0800 ;
        RECT 5.8150 1.8000 5.9150 2.0800 ;
        RECT 6.1200 1.8000 6.2200 2.0800 ;
        RECT 6.6400 1.8000 6.7400 2.0800 ;
        RECT 0.0750 1.7900 0.1750 2.0800 ;
        RECT 0.5950 1.7900 0.6950 2.0800 ;
        RECT 1.1150 1.7900 1.2150 2.0800 ;
        RECT 1.6350 1.7900 1.7350 2.0800 ;
        RECT 2.1550 1.7900 2.2550 2.0800 ;
        RECT 2.6750 1.7900 2.7750 2.0800 ;
        RECT 3.1950 1.7900 3.2950 2.0800 ;
        RECT 7.1850 1.7550 7.2850 2.0800 ;
        RECT 7.7050 1.7550 7.8050 2.0800 ;
        RECT 8.2250 1.7350 8.3250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2550 0.9750 0.3450 1.2150 ;
      RECT 0.2550 0.8850 4.2000 0.9750 ;
      RECT 4.1100 0.8200 4.2000 0.8850 ;
      RECT 4.1100 1.4400 5.6900 1.5300 ;
      RECT 4.1100 0.7300 5.7500 0.8200 ;
      RECT 4.1100 0.9750 4.2000 1.4400 ;
      RECT 4.7400 0.4100 4.8300 0.7300 ;
      RECT 5.6600 0.4100 5.7500 0.7300 ;
      RECT 0.9850 0.8850 1.3550 1.1350 ;
      RECT 2.0250 0.8850 2.3950 1.1350 ;
      RECT 3.0650 0.8850 3.4350 1.1350 ;
      RECT 0.4450 1.0950 0.8550 1.1850 ;
      RECT 0.7650 1.2250 3.9550 1.3150 ;
      RECT 0.7650 1.1850 0.8550 1.2250 ;
      RECT 3.8650 1.6600 7.0200 1.7100 ;
      RECT 3.8650 1.6200 8.0600 1.6600 ;
      RECT 3.8650 1.3150 3.9550 1.6200 ;
      RECT 6.9300 1.7100 7.0200 1.9600 ;
      RECT 6.9300 0.8400 7.0200 1.5700 ;
      RECT 6.9300 1.5700 8.0600 1.6200 ;
      RECT 6.9300 0.7500 7.5400 0.8400 ;
      RECT 7.4500 1.2000 8.0400 1.2900 ;
      RECT 7.4500 1.6600 7.5400 1.9800 ;
      RECT 7.4500 0.8400 7.5400 1.2000 ;
      RECT 7.9500 0.8400 8.0400 1.2000 ;
      RECT 7.9500 0.7500 8.3200 0.8400 ;
      RECT 7.9700 1.6600 8.0600 1.9800 ;
      RECT 1.5050 1.0950 1.8750 1.3150 ;
      RECT 2.5450 1.0950 2.9150 1.3150 ;
      RECT 3.5850 1.0950 3.9550 1.3150 ;
      RECT 8.4400 0.9700 8.7250 1.0650 ;
      RECT 6.7500 0.5600 8.5300 0.6500 ;
      RECT 8.4400 0.6500 8.5300 0.9700 ;
      RECT 6.3000 1.3700 6.8400 1.4600 ;
      RECT 6.7450 0.9300 6.8400 1.3700 ;
      RECT 6.3850 0.8400 6.8400 0.9300 ;
      RECT 6.7500 0.6500 6.8400 0.8400 ;
      RECT 6.3850 0.4750 6.4750 0.8400 ;
      RECT 7.7700 0.6500 7.8600 1.0100 ;
      RECT 7.6500 1.0100 7.8600 1.1100 ;
  END
END MX2_X8B_A12TH

MACRO MXIT2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7550 ;
        RECT 1.8050 0.3200 1.9050 0.8550 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0650 0.5800 1.4000 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END B

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9550 0.3500 1.2550 ;
        RECT 0.2500 0.8650 0.6300 0.9550 ;
        RECT 0.5400 0.5700 0.6300 0.8650 ;
        RECT 0.5400 0.4800 1.0300 0.5700 ;
        RECT 0.9400 0.5700 1.0300 0.9950 ;
        RECT 0.9400 0.9950 1.2700 1.0850 ;
        RECT 1.1800 1.0850 1.2700 1.5100 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1400 1.6200 1.4600 1.7500 ;
        RECT 1.1400 1.7500 1.2300 1.9900 ;
        RECT 1.3600 0.7500 1.4600 1.6200 ;
        RECT 1.1350 0.6500 1.4600 0.7500 ;
    END
    ANTENNADIFFAREA 0.1782 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1800 1.9500 1.4200 ;
        RECT 1.7300 1.0800 1.9500 1.1800 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.8050 1.5750 1.9050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7400 0.6700 0.8300 1.6950 ;
      RECT 0.0550 1.7850 1.0400 1.8750 ;
      RECT 0.9500 1.1950 1.0400 1.7850 ;
      RECT 0.0550 0.7550 0.1450 1.7850 ;
      RECT 0.0550 0.6650 0.2450 0.7550 ;
      RECT 1.5500 0.4450 1.6400 1.9600 ;
  END
END MXIT2_X0P5M_A12TH

MACRO LATRPQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7800 ;
        RECT 0.6750 0.3200 0.7650 0.6000 ;
        RECT 1.1950 0.3200 1.2850 0.6000 ;
        RECT 2.4350 0.3200 2.5350 0.8400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 2.3900 2.0250 2.6000 2.0800 ;
        RECT 0.6200 1.8950 0.7900 2.0800 ;
        RECT 1.1950 1.7950 1.2850 2.0800 ;
    END
  END VDD

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2200 0.5500 1.3950 ;
        RECT 0.4500 1.0500 0.6050 1.2200 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.1500 2.5500 1.6250 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.8100 2.1500 1.2300 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7800 1.3500 1.4350 ;
        RECT 0.8750 1.4350 1.3500 1.5250 ;
        RECT 0.9350 0.6900 1.3500 0.7800 ;
        RECT 0.9350 0.4100 1.0250 0.6900 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN
  OBS
    LAYER M1 ;
      RECT 0.0550 0.8700 0.9500 0.9600 ;
      RECT 0.8600 0.9600 0.9500 1.1600 ;
      RECT 0.0550 1.6050 0.1700 1.9750 ;
      RECT 0.0550 0.9600 0.1450 1.6050 ;
      RECT 0.3400 0.5300 0.4300 0.8700 ;
      RECT 0.2600 1.7000 1.5300 1.7050 ;
      RECT 0.9700 1.6500 1.5300 1.7000 ;
      RECT 0.9700 1.6150 1.9200 1.6500 ;
      RECT 1.8300 1.6500 1.9200 1.9650 ;
      RECT 1.4400 1.5600 1.9200 1.6150 ;
      RECT 1.4400 0.7500 1.5300 1.5600 ;
      RECT 1.4400 0.6600 1.9450 0.7500 ;
      RECT 1.8550 0.7500 1.9450 0.8300 ;
      RECT 1.8550 0.4150 1.9450 0.6600 ;
      RECT 0.2600 1.0700 0.3500 1.7000 ;
      RECT 0.2600 1.7050 1.0600 1.7900 ;
      RECT 2.1900 1.4400 2.2800 1.7200 ;
      RECT 2.1900 1.3500 2.3300 1.4400 ;
      RECT 2.2400 0.6750 2.3300 1.3500 ;
      RECT 2.0650 0.5850 2.3300 0.6750 ;
      RECT 2.0100 1.8300 2.9500 1.9200 ;
      RECT 2.8300 1.7150 2.9500 1.8300 ;
      RECT 2.8600 0.7550 2.9500 1.7150 ;
      RECT 2.8300 0.5650 2.9500 0.7550 ;
      RECT 2.0100 1.4500 2.1000 1.8300 ;
      RECT 1.6500 1.3600 2.1000 1.4500 ;
      RECT 1.6500 0.8600 1.7400 1.3600 ;
  END
END LATRPQN_X2M_A12TH

MACRO LATRPQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6950 ;
        RECT 0.8600 0.3200 0.9500 0.6000 ;
        RECT 1.3950 0.3200 1.4850 0.4450 ;
        RECT 1.6250 0.3200 1.7150 0.6750 ;
        RECT 2.7300 0.3200 2.8200 0.9000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3400 1.8400 0.4300 2.0800 ;
        RECT 0.8600 1.7550 0.9500 2.0800 ;
        RECT 1.5900 1.5400 1.6800 2.0800 ;
    END
  END VDD

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.6900 0.9500 1.0350 ;
        RECT 0.8500 1.0350 1.0250 1.2050 ;
    END
    ANTENNAGATEAREA 0.0774 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.2100 2.7500 1.6300 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 0.8050 2.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.6500 0.7300 1.7500 ;
        RECT 0.5600 1.7500 0.7300 1.9400 ;
        RECT 0.0800 1.0000 0.1700 1.6500 ;
        RECT 0.0800 0.9100 0.6900 1.0000 ;
        RECT 0.0800 0.5300 0.1700 0.9100 ;
        RECT 0.6000 0.5300 0.6900 0.9100 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN
  OBS
    LAYER M1 ;
      RECT 1.2550 0.7700 1.7000 0.8600 ;
      RECT 0.6100 1.1800 0.7000 1.4700 ;
      RECT 0.3100 1.0900 0.7000 1.1800 ;
      RECT 1.3300 1.5600 1.4200 1.7350 ;
      RECT 0.6100 1.4700 1.4200 1.5600 ;
      RECT 1.2550 1.2800 1.4200 1.4700 ;
      RECT 1.2550 0.8600 1.3450 1.2800 ;
      RECT 1.2550 0.6200 1.3450 0.7700 ;
      RECT 1.0750 0.5300 1.3450 0.6200 ;
      RECT 1.8250 0.5150 2.2400 0.6050 ;
      RECT 2.1100 1.6400 2.2000 1.9600 ;
      RECT 1.8250 1.5500 2.2000 1.6400 ;
      RECT 1.8250 1.1100 1.9150 1.5500 ;
      RECT 1.4350 1.0200 1.9150 1.1100 ;
      RECT 1.8250 0.6050 1.9150 1.0200 ;
      RECT 2.4700 1.1550 2.5600 1.7150 ;
      RECT 2.4400 1.0650 2.5600 1.1550 ;
      RECT 2.4400 0.7000 2.5300 1.0650 ;
      RECT 3.0300 1.9150 3.1500 1.9900 ;
      RECT 2.2900 1.8250 3.1500 1.9150 ;
      RECT 3.0300 1.5700 3.1500 1.8250 ;
      RECT 3.0600 0.9250 3.1500 1.5700 ;
      RECT 3.0300 0.5350 3.1500 0.9250 ;
      RECT 2.2900 1.4500 2.3800 1.8250 ;
      RECT 2.0250 1.3600 2.3800 1.4500 ;
      RECT 2.0250 0.7250 2.1150 1.3600 ;
  END
END LATRPQN_X3M_A12TH

MACRO LATRPQN_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.3600 ;
        RECT 1.5550 0.3200 1.6450 0.6400 ;
        RECT 1.8100 0.3200 1.9000 0.6200 ;
        RECT 2.3300 0.3200 2.4200 0.6200 ;
        RECT 2.5900 0.3200 2.6800 0.6350 ;
        RECT 3.1100 0.3200 3.2000 0.6550 ;
        RECT 3.6300 0.3200 3.7200 0.6550 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8500 0.5900 0.9500 ;
        RECT 0.2500 0.7200 0.3400 0.8500 ;
    END
    ANTENNAGATEAREA 0.1014 ;
  END G

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.1500 0.3500 1.3900 ;
        RECT 0.2500 1.0500 0.5900 1.1500 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0900 2.5550 1.1900 ;
        RECT 2.4650 1.0200 2.5550 1.0900 ;
        RECT 1.8500 0.9500 1.9650 1.0900 ;
    END
    ANTENNAGATEAREA 0.1272 ;
  END R

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.2500 3.5850 1.3500 ;
        RECT 2.8500 1.3500 2.9400 1.7450 ;
        RECT 3.3700 1.3500 3.4600 1.7550 ;
        RECT 3.4950 0.9800 3.5850 1.2500 ;
        RECT 2.8500 0.8900 3.5850 0.9800 ;
        RECT 2.8500 0.5200 2.9400 0.8900 ;
        RECT 3.3700 0.5200 3.4600 0.8900 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.3800 1.8950 0.5500 2.0800 ;
        RECT 2.5900 1.7750 2.6800 2.0800 ;
        RECT 3.1100 1.7650 3.2000 2.0800 ;
        RECT 3.6300 1.7650 3.7200 2.0800 ;
        RECT 1.6350 1.6100 1.7250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6450 1.3350 0.8150 1.6250 ;
      RECT 0.7250 0.8100 0.8150 1.3350 ;
      RECT 0.6850 0.4400 0.8150 0.8100 ;
      RECT 0.0500 1.7150 1.0150 1.8050 ;
      RECT 0.9250 1.4800 1.0150 1.7150 ;
      RECT 0.9250 1.3900 1.1950 1.4800 ;
      RECT 1.1050 0.8850 1.1950 1.3900 ;
      RECT 0.0500 1.8050 0.1700 1.9300 ;
      RECT 0.0500 1.5600 0.1700 1.7150 ;
      RECT 0.0500 0.6500 0.1500 1.5600 ;
      RECT 0.0500 0.4400 0.1700 0.6500 ;
      RECT 1.3300 1.2800 2.2600 1.3700 ;
      RECT 1.1050 1.6600 1.1950 1.9900 ;
      RECT 1.1050 1.5700 1.4200 1.6600 ;
      RECT 1.3300 1.3700 1.4200 1.5700 ;
      RECT 1.3300 0.7800 1.4200 1.2800 ;
      RECT 0.9050 0.6900 1.4200 0.7800 ;
      RECT 2.6650 1.0700 3.3850 1.1600 ;
      RECT 1.5200 0.8200 1.6100 1.0900 ;
      RECT 2.1100 1.6650 2.2000 1.9800 ;
      RECT 2.0700 0.4100 2.1600 0.7300 ;
      RECT 2.1100 1.5750 2.7550 1.6650 ;
      RECT 2.6650 1.1600 2.7550 1.5750 ;
      RECT 2.6650 0.8200 2.7550 1.0700 ;
      RECT 1.5200 0.7300 2.7550 0.8200 ;
  END
END LATRPQN_X4M_A12TH

MACRO LATRQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.7050 0.3200 0.7950 0.3900 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7150 0.1500 1.5800 ;
        RECT 0.0500 1.5800 0.1750 1.9700 ;
        RECT 0.0500 0.5050 0.1750 0.7150 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2350 0.9900 2.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8900 2.7650 0.9900 ;
        RECT 2.4500 0.5800 2.5500 0.8900 ;
        RECT 2.6700 0.9900 2.7650 1.3000 ;
        RECT 1.7800 0.4800 2.5500 0.5800 ;
        RECT 1.7800 0.5800 1.8700 0.6400 ;
        RECT 1.5400 0.6400 1.8700 0.7300 ;
        RECT 1.5400 0.7300 1.6400 0.9950 ;
        RECT 0.8600 0.9950 1.6400 1.0950 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END G

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.2500 1.6950 1.3600 ;
        RECT 1.6050 1.3600 1.6950 1.6350 ;
        RECT 0.7000 1.2350 0.8700 1.2500 ;
        RECT 1.6050 1.6350 2.5750 1.7250 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END RN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 1.2000 1.8400 1.3000 2.0800 ;
        RECT 2.1100 1.8400 2.2000 2.0800 ;
        RECT 2.5700 1.8300 2.6600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5200 0.6600 1.1800 0.7500 ;
      RECT 1.0900 0.7500 1.1800 0.8950 ;
      RECT 0.5200 1.6300 0.7850 1.7200 ;
      RECT 0.5200 0.7500 0.6100 1.6300 ;
      RECT 0.3400 0.4800 1.6700 0.5000 ;
      RECT 1.4050 1.8350 1.6150 1.9250 ;
      RECT 1.3550 0.4100 1.6700 0.4800 ;
      RECT 0.9950 1.5850 1.4950 1.6750 ;
      RECT 0.3400 0.5000 1.4450 0.5700 ;
      RECT 1.4050 1.6750 1.4950 1.8350 ;
      RECT 0.3400 0.5700 0.4300 1.8300 ;
      RECT 0.6450 1.9200 0.8150 1.9750 ;
      RECT 0.3400 1.8300 1.0850 1.9200 ;
      RECT 0.9950 1.6750 1.0850 1.8300 ;
      RECT 1.8050 0.9100 1.8950 1.5450 ;
      RECT 1.8050 0.8200 2.0500 0.9100 ;
      RECT 1.9600 0.6900 2.0500 0.8200 ;
      RECT 2.8300 1.8850 2.9200 1.9900 ;
      RECT 2.8300 1.7950 2.9550 1.8850 ;
      RECT 2.8650 1.5400 2.9550 1.7950 ;
      RECT 2.0050 1.4500 2.9550 1.5400 ;
      RECT 2.8650 0.6000 2.9550 1.4500 ;
      RECT 2.8300 0.4300 2.9550 0.6000 ;
      RECT 2.0050 1.0600 2.0950 1.4500 ;
  END
END LATRQ_X0P5M_A12TH

MACRO LATRQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.3900 ;
        RECT 0.7050 0.3200 0.7950 0.3900 ;
        RECT 2.5800 0.3200 2.6700 0.3900 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9150 0.1500 1.2900 ;
        RECT 0.0500 1.2900 0.1750 1.7200 ;
        RECT 0.0500 0.4850 0.1750 0.9150 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2450 0.9000 2.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.5800 2.5500 0.9450 ;
        RECT 2.4500 0.9450 2.7650 1.0450 ;
        RECT 1.8300 0.4800 2.5500 0.5800 ;
        RECT 2.6700 1.0450 2.7650 1.3350 ;
        RECT 1.8300 0.5800 1.9200 0.6100 ;
        RECT 1.5850 0.6100 1.9200 0.7000 ;
        RECT 1.5850 0.7000 1.6850 0.9950 ;
        RECT 0.8600 0.9950 1.6850 1.0950 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END G

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.2500 1.6950 1.3600 ;
        RECT 1.6050 1.3600 1.6950 1.6350 ;
        RECT 0.7000 1.2350 0.8700 1.2500 ;
        RECT 1.6050 1.6350 2.5750 1.7250 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END RN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.3350 1.9450 0.4350 2.0800 ;
        RECT 2.0650 1.8400 2.1550 2.0800 ;
        RECT 2.5700 1.8150 2.6600 2.0800 ;
        RECT 1.2000 1.7650 1.3000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5200 0.6600 1.1800 0.7500 ;
      RECT 1.0900 0.7500 1.1800 0.8950 ;
      RECT 0.5200 1.4950 0.7850 1.5850 ;
      RECT 0.5200 0.7500 0.6100 1.4950 ;
      RECT 1.4250 1.8350 1.6150 1.9250 ;
      RECT 0.3400 0.4800 1.7100 0.5200 ;
      RECT 1.3700 0.4300 1.7100 0.4800 ;
      RECT 1.4250 1.6750 1.5150 1.8350 ;
      RECT 0.9950 1.5850 1.5150 1.6750 ;
      RECT 0.3400 0.5200 1.4600 0.5700 ;
      RECT 0.3400 0.5700 0.4300 1.7350 ;
      RECT 0.6850 1.8250 0.7750 1.9750 ;
      RECT 0.9950 1.6750 1.0850 1.7350 ;
      RECT 0.3400 1.7350 1.0850 1.8250 ;
      RECT 1.8050 0.8800 1.8950 1.5450 ;
      RECT 1.8050 0.7900 2.1000 0.8800 ;
      RECT 2.0100 0.6900 2.1000 0.7900 ;
      RECT 2.8300 1.8850 2.9200 1.9900 ;
      RECT 2.8300 1.7950 2.9550 1.8850 ;
      RECT 2.8650 1.5400 2.9550 1.7950 ;
      RECT 2.0050 1.4500 2.9550 1.5400 ;
      RECT 2.8650 0.8600 2.9550 1.4500 ;
      RECT 2.8300 0.6350 2.9550 0.8600 ;
      RECT 2.0050 0.9700 2.0950 1.4500 ;
  END
END LATRQ_X1M_A12TH

MACRO LATRQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4400 0.4200 ;
        RECT 2.0200 0.3200 2.1200 0.4200 ;
        RECT 2.4100 0.3200 2.5800 0.3600 ;
        RECT 2.9700 0.3200 3.0600 0.6900 ;
    END
  END VSS

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0250 0.5500 1.4500 ;
        RECT 0.4500 1.4500 0.7300 1.5500 ;
        RECT 0.6300 1.5500 0.7300 1.6200 ;
        RECT 0.6300 1.6200 1.9750 1.7200 ;
        RECT 1.8850 1.7200 1.9750 1.9400 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END RN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9050 0.7700 1.2550 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7100 1.0500 2.9950 1.1500 ;
        RECT 2.7100 1.1500 2.8000 1.7200 ;
        RECT 2.7100 0.5500 2.8000 1.0500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.6100 0.3500 1.8200 ;
        RECT 0.0900 1.8200 1.4450 1.9200 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3600 2.0400 0.7700 2.0800 ;
        RECT 1.6050 1.8450 1.7750 2.0800 ;
        RECT 2.4500 1.7900 2.5400 2.0800 ;
        RECT 2.9700 1.7700 3.0600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8400 1.4400 1.0100 1.5300 ;
      RECT 0.8600 0.9200 0.9500 1.4400 ;
      RECT 0.8600 0.7100 0.9700 0.9200 ;
      RECT 1.0400 1.2100 1.2150 1.3000 ;
      RECT 1.0800 0.5700 1.1700 1.2100 ;
      RECT 0.6500 0.4800 1.5800 0.5700 ;
      RECT 0.6500 0.5700 0.7400 0.6100 ;
      RECT 1.4900 0.5700 1.5800 0.8300 ;
      RECT 0.0950 0.6100 0.7400 0.7000 ;
      RECT 0.0950 0.7000 0.1850 1.5100 ;
      RECT 1.1500 1.4400 2.0600 1.5300 ;
      RECT 1.9700 1.1700 2.0600 1.4400 ;
      RECT 1.3400 1.0000 1.4300 1.4400 ;
      RECT 1.9700 1.0800 2.3750 1.1700 ;
      RECT 1.2600 0.9100 1.4300 1.0000 ;
      RECT 1.2600 0.7100 1.3500 0.9100 ;
      RECT 2.1500 1.3200 2.5750 1.4100 ;
      RECT 2.4850 0.9400 2.5750 1.3200 ;
      RECT 1.7200 0.8500 2.5750 0.9400 ;
      RECT 1.7200 0.9400 1.8100 0.9500 ;
      RECT 1.5350 0.9500 1.8100 1.0400 ;
      RECT 1.5350 1.0400 1.6250 1.1300 ;
  END
END LATRQ_X2M_A12TH

MACRO LATRQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4400 0.4200 ;
        RECT 2.0200 0.3200 2.1200 0.4200 ;
        RECT 2.4100 0.3200 2.5800 0.3600 ;
        RECT 2.9700 0.3200 3.0600 0.6850 ;
    END
  END VSS

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0250 0.5500 1.4500 ;
        RECT 0.4500 1.4500 0.7300 1.5500 ;
        RECT 0.6300 1.5500 0.7300 1.6200 ;
        RECT 0.6300 1.6200 1.9750 1.7200 ;
        RECT 1.8850 1.7200 1.9750 1.9400 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END RN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9050 0.7700 1.2550 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7100 1.0500 3.3200 1.1500 ;
        RECT 2.7100 1.1500 2.8000 1.7200 ;
        RECT 3.2300 1.1500 3.3200 1.7200 ;
        RECT 2.7100 0.5400 2.8000 1.0500 ;
        RECT 3.2300 0.5400 3.3200 1.0500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.6100 0.3500 1.8200 ;
        RECT 0.0900 1.8200 1.4450 1.9200 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.6050 1.8450 1.7750 2.0800 ;
        RECT 2.4500 1.7900 2.5400 2.0800 ;
        RECT 2.9700 1.7700 3.0600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8400 1.4400 1.0300 1.5300 ;
      RECT 0.8600 0.9400 0.9500 1.4400 ;
      RECT 0.8600 0.7300 0.9700 0.9400 ;
      RECT 1.0400 1.2100 1.2350 1.3000 ;
      RECT 1.0600 0.5700 1.1500 1.2100 ;
      RECT 0.6500 0.4800 1.5800 0.5700 ;
      RECT 0.6500 0.5700 0.7400 0.5950 ;
      RECT 1.4900 0.5700 1.5800 0.8300 ;
      RECT 0.0950 0.5950 0.7400 0.6850 ;
      RECT 0.0950 0.6850 0.1850 1.5100 ;
      RECT 1.1400 1.4400 2.0600 1.5300 ;
      RECT 1.9700 1.1700 2.0600 1.4400 ;
      RECT 1.3400 1.0000 1.4300 1.4400 ;
      RECT 1.9700 1.0800 2.3750 1.1700 ;
      RECT 1.2600 0.9100 1.4300 1.0000 ;
      RECT 1.2600 0.7300 1.3500 0.9100 ;
      RECT 2.1500 1.3200 2.5750 1.4100 ;
      RECT 2.4850 0.9400 2.5750 1.3200 ;
      RECT 1.7200 0.8500 2.5750 0.9400 ;
      RECT 1.7200 0.9400 1.8100 0.9500 ;
      RECT 1.5350 0.9500 1.8100 1.0400 ;
      RECT 1.5350 1.0400 1.6250 1.3300 ;
  END
END LATRQ_X3M_A12TH

MACRO LATSPQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 1.8300 0.3200 2.0000 0.4550 ;
        RECT 2.4800 0.3200 2.6500 0.7550 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.8500 1.4000 1.9500 ;
        RECT 1.0100 1.8100 1.1100 1.8500 ;
        RECT 0.1150 1.7100 1.1100 1.8100 ;
        RECT 0.1150 1.5600 0.2850 1.7100 ;
    END
    ANTENNAGATEAREA 0.0417 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.3100 1.9000 0.4800 2.0800 ;
        RECT 2.5150 1.5350 2.6150 2.0800 ;
        RECT 1.9500 1.5100 2.0500 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0050 2.9500 1.2550 ;
        RECT 2.7750 1.2550 2.9500 1.3550 ;
        RECT 2.7750 0.9050 2.9500 1.0050 ;
        RECT 2.7750 1.3550 2.8750 1.7300 ;
        RECT 2.7750 0.5750 2.8750 0.9050 ;
    END
    ANTENNADIFFAREA 0.14175 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 0.8500 0.7250 1.0000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3300 1.6500 1.8600 1.7500 ;
        RECT 1.3300 1.6200 1.4200 1.6500 ;
        RECT 0.4450 1.5200 1.4200 1.6200 ;
        RECT 0.4450 1.0900 0.5450 1.5200 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END S
  OBS
    LAYER M1 ;
      RECT 0.8150 1.3400 0.9950 1.4300 ;
      RECT 0.8150 0.8500 0.9050 1.3400 ;
      RECT 0.8150 0.6800 0.9550 0.8500 ;
      RECT 0.0800 0.4800 1.5900 0.5700 ;
      RECT 1.0500 0.5700 1.1400 1.2300 ;
      RECT 1.5000 0.5700 1.5900 0.7400 ;
      RECT 0.0800 0.5700 0.1700 1.4600 ;
      RECT 1.9650 1.0800 2.5000 1.1700 ;
      RECT 1.1050 1.3400 1.3250 1.4300 ;
      RECT 1.2350 0.9250 1.3250 1.3400 ;
      RECT 1.2350 0.6800 1.3250 0.8350 ;
      RECT 1.2350 0.8350 2.0550 0.9250 ;
      RECT 1.9650 0.9250 2.0550 1.0800 ;
      RECT 1.9650 0.6550 2.0550 0.8350 ;
      RECT 1.9650 0.5650 2.2700 0.6550 ;
      RECT 2.1000 0.4200 2.2700 0.5650 ;
      RECT 1.5250 1.3200 2.6850 1.4100 ;
      RECT 1.5250 1.0150 1.6150 1.3200 ;
      RECT 2.5950 0.9400 2.6850 1.3200 ;
      RECT 2.1450 0.8500 2.6850 0.9400 ;
  END
END LATSPQ_X0P5M_A12TH

MACRO LATSPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
    END
  END VSS

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5800 0.1600 1.3000 ;
        RECT 0.0500 0.5100 0.8450 0.5800 ;
        RECT 0.0500 0.4800 1.1250 0.5100 ;
        RECT 0.7550 0.4100 1.1250 0.4800 ;
    END
    ANTENNAGATEAREA 0.0786 ;
  END S

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0800 0.3500 1.3000 ;
        RECT 0.2500 0.8950 0.4450 1.0800 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9150 3.1500 1.2900 ;
        RECT 2.9950 1.2900 3.1500 1.4400 ;
        RECT 2.9950 0.7650 3.1500 0.9150 ;
        RECT 2.9950 1.4400 3.0950 1.7200 ;
        RECT 2.9950 0.4850 3.0950 0.7650 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Q

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9000 1.9650 1.3000 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.6350 1.8500 1.8050 2.0800 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 2.7350 1.7700 2.8350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5400 0.7600 0.6300 1.6750 ;
      RECT 0.3650 0.6700 0.6300 0.7600 ;
      RECT 1.1250 1.2950 1.5300 1.3850 ;
      RECT 1.1250 0.9750 1.2150 1.2950 ;
      RECT 1.0450 0.8850 1.2150 0.9750 ;
      RECT 0.9800 1.4800 2.2200 1.5700 ;
      RECT 2.1300 0.6700 2.2200 1.4800 ;
      RECT 1.6450 1.0300 1.7350 1.4800 ;
      RECT 0.6350 1.8000 1.0700 1.8900 ;
      RECT 0.9800 1.5700 1.0700 1.8000 ;
      RECT 1.1650 1.6600 2.4650 1.7500 ;
      RECT 2.3750 0.7350 2.4650 1.6600 ;
      RECT 1.1650 1.7500 1.3350 1.8550 ;
      RECT 2.5550 1.0800 2.9450 1.1700 ;
      RECT 2.5550 0.5700 2.6450 1.0800 ;
      RECT 1.7900 0.4800 2.6450 0.5700 ;
      RECT 1.7900 0.5700 1.8800 0.6700 ;
      RECT 0.8000 0.6700 1.8800 0.7600 ;
      RECT 0.8000 0.7600 0.8900 1.6350 ;
  END
END LATSPQ_X1M_A12TH

MACRO LATSPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 1.8050 0.3200 2.0150 0.5300 ;
        RECT 2.4900 0.3200 2.5900 0.6750 ;
        RECT 3.0100 0.3200 3.1100 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.4900 1.7700 2.5900 2.0800 ;
        RECT 3.0100 1.7700 3.1100 2.0800 ;
        RECT 1.9350 1.5000 2.0350 2.0800 ;
    END
  END VDD

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.6100 1.8400 1.7100 ;
        RECT 1.5800 1.7100 1.8400 1.7500 ;
        RECT 0.4500 1.0500 0.5500 1.6100 ;
    END
    ANTENNAGATEAREA 0.0786 ;
  END S

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7600 0.7500 1.1800 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9800 2.9500 1.2600 ;
        RECT 2.7500 1.2600 2.9500 1.3600 ;
        RECT 2.7500 0.8800 2.9500 0.9800 ;
        RECT 2.7500 1.3600 2.8500 1.7300 ;
        RECT 2.7500 0.5400 2.8500 0.8800 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1950 1.8100 1.4000 1.9100 ;
        RECT 0.1950 1.9100 0.5950 1.9500 ;
        RECT 0.1950 1.7250 0.2950 1.8100 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END G
  OBS
    LAYER M1 ;
      RECT 0.8600 0.6650 0.9500 1.5000 ;
      RECT 1.4600 0.6900 1.6500 0.7800 ;
      RECT 1.4600 0.5700 1.5500 0.6900 ;
      RECT 0.0950 0.5600 1.5500 0.5700 ;
      RECT 0.0950 0.5700 0.7400 0.6500 ;
      RECT 1.0600 0.5700 1.1500 1.2300 ;
      RECT 0.6500 0.4800 1.5500 0.5600 ;
      RECT 0.0950 0.6500 0.1850 1.6350 ;
      RECT 1.2600 0.8900 1.9650 0.9800 ;
      RECT 1.8750 0.9800 1.9650 1.0800 ;
      RECT 1.8750 0.7350 1.9650 0.8900 ;
      RECT 1.8750 1.0800 2.4550 1.1700 ;
      RECT 1.8750 0.6450 2.2250 0.7350 ;
      RECT 2.1350 0.4100 2.2250 0.6450 ;
      RECT 1.1000 1.3700 1.3500 1.4600 ;
      RECT 1.2600 0.9800 1.3500 1.3700 ;
      RECT 1.2600 0.6650 1.3500 0.8900 ;
      RECT 1.5300 1.3200 2.6550 1.4100 ;
      RECT 1.5300 1.0700 1.6200 1.3200 ;
      RECT 2.5650 0.9400 2.6550 1.3200 ;
      RECT 2.0950 0.8500 2.6550 0.9400 ;
  END
END LATSPQ_X2M_A12TH

MACRO LATSPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.4300 0.3200 0.5950 0.4650 ;
        RECT 1.0400 0.3200 1.2100 0.4650 ;
        RECT 2.3150 0.3200 2.4150 0.8000 ;
        RECT 3.2300 0.3200 3.3300 0.6850 ;
        RECT 3.7500 0.3200 3.8500 0.6900 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4900 1.2500 4.1500 1.3500 ;
        RECT 3.4900 1.3500 3.5900 1.7350 ;
        RECT 4.0100 1.3500 4.1500 1.7450 ;
        RECT 3.4900 0.5900 3.5900 1.2500 ;
        RECT 4.0100 0.5900 4.1500 1.2500 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 3.2300 1.7650 3.3350 2.0800 ;
        RECT 3.7500 1.7650 3.8500 2.0800 ;
        RECT 2.6400 1.5000 2.8100 2.0800 ;
    END
  END VDD

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.6000 2.5500 1.9300 ;
        RECT 0.4400 1.5000 2.5500 1.6000 ;
        RECT 0.4400 0.9900 0.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.1332 ;
  END S

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.0500 1.1400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1400 1.8500 0.4600 1.9500 ;
        RECT 0.3650 1.7500 1.9050 1.8500 ;
        RECT 1.8050 1.8500 2.2200 1.9500 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END G
  OBS
    LAYER M1 ;
      RECT 0.0950 0.5550 1.5750 0.6450 ;
      RECT 1.4850 0.5400 1.5750 0.5550 ;
      RECT 1.4850 0.4500 1.9000 0.5400 ;
      RECT 0.0950 0.6450 0.1850 1.7200 ;
      RECT 1.6650 0.8900 2.7150 0.9800 ;
      RECT 2.6250 0.9800 2.7150 1.0800 ;
      RECT 2.6250 0.6450 2.7150 0.8900 ;
      RECT 2.6250 1.0800 3.2150 1.1700 ;
      RECT 1.8950 1.3000 2.0850 1.4100 ;
      RECT 1.9950 0.9800 2.0850 1.3000 ;
      RECT 1.6650 0.6750 1.7550 0.8900 ;
      RECT 2.2900 1.3200 3.4000 1.4100 ;
      RECT 2.2900 1.0700 2.3800 1.3200 ;
      RECT 3.3100 0.9400 3.4000 1.3200 ;
      RECT 2.8250 0.8500 3.4000 0.9400 ;
      RECT 0.7400 1.3200 1.7950 1.4100 ;
      RECT 1.3350 1.3000 1.7950 1.3200 ;
      RECT 1.3350 0.8850 1.4400 1.3000 ;
      RECT 0.7350 0.7950 1.4400 0.8850 ;
  END
END LATSPQ_X3M_A12TH

MACRO LATSQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 1.1400 0.3200 1.2300 0.6500 ;
        RECT 0.3400 0.3200 0.4300 0.5200 ;
        RECT 2.2950 0.3200 2.3850 0.7500 ;
        RECT 0.8850 0.6500 1.2300 0.7400 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.3400 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 1.2500 2.4300 1.3500 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0950 0.8500 2.5400 0.9500 ;
        RECT 2.4500 0.9500 2.5400 1.1000 ;
        RECT 2.0950 0.5700 2.1850 0.8500 ;
        RECT 1.6300 0.4800 2.1850 0.5700 ;
        RECT 1.6300 0.5700 1.7300 1.0800 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.4200 0.1700 1.9200 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.3000 1.7150 2.3900 2.0800 ;
        RECT 0.3400 1.7050 0.4300 2.0800 ;
        RECT 0.9200 1.5950 1.0300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6600 0.8800 1.0400 0.9700 ;
      RECT 0.6600 0.4200 1.0300 0.5100 ;
      RECT 0.6000 1.9000 0.8100 1.9900 ;
      RECT 0.6600 1.5600 0.7500 1.9000 ;
      RECT 0.3000 1.4700 0.7500 1.5600 ;
      RECT 0.6600 0.9700 0.7500 1.4700 ;
      RECT 0.6600 0.5100 0.7500 0.8800 ;
      RECT 1.4250 1.4900 1.5150 1.7900 ;
      RECT 1.1500 1.4000 1.5150 1.4900 ;
      RECT 1.1500 1.1500 1.2400 1.4000 ;
      RECT 0.8450 1.0600 1.2400 1.1500 ;
      RECT 1.1500 0.9250 1.2400 1.0600 ;
      RECT 1.1500 0.8350 1.5200 0.9250 ;
      RECT 1.4300 0.6200 1.5200 0.8350 ;
      RECT 0.8450 1.1500 0.9350 1.2600 ;
      RECT 1.8300 1.6400 2.0100 1.7300 ;
      RECT 1.8300 0.7700 1.9200 1.6400 ;
      RECT 1.8300 0.6800 2.0000 0.7700 ;
      RECT 2.1200 1.5150 2.7200 1.6050 ;
      RECT 2.6300 1.6050 2.7200 1.8150 ;
      RECT 2.6300 0.6050 2.7200 1.5150 ;
      RECT 1.3700 1.0150 1.4600 1.1900 ;
      RECT 1.6500 1.2800 1.7400 1.8200 ;
      RECT 1.3700 1.1900 1.7400 1.2800 ;
      RECT 1.6500 1.8200 2.2100 1.9100 ;
      RECT 2.1200 1.6050 2.2100 1.8200 ;
  END
END LATSQN_X0P5M_A12TH

MACRO LATSQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3450 0.3200 0.4350 0.6350 ;
        RECT 1.0450 0.3200 1.1350 0.6900 ;
        RECT 2.3500 0.3200 2.4400 0.7200 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.5600 1.3450 ;
    END
    ANTENNAGATEAREA 0.0558 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1250 1.2500 2.5300 1.3500 ;
        RECT 2.1250 1.0950 2.2150 1.2500 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8100 1.8250 0.9950 ;
        RECT 1.7350 0.5700 1.8250 0.8100 ;
        RECT 1.7350 0.4800 2.2400 0.5700 ;
        RECT 2.1500 0.5700 2.2400 0.8500 ;
        RECT 2.1500 0.8500 2.5500 0.9500 ;
        RECT 2.4450 0.9500 2.5500 1.0950 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9100 0.1500 1.6500 ;
        RECT 0.0500 1.6500 0.1950 1.9900 ;
        RECT 0.0500 0.4950 0.1750 0.9100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.3050 1.7000 2.3950 2.0800 ;
        RECT 0.3450 1.6850 0.4350 2.0800 ;
        RECT 0.8850 1.5350 0.9750 2.0800 ;
        RECT 0.8850 1.4200 1.1350 1.5350 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6750 0.9000 1.1350 0.9900 ;
      RECT 1.0450 0.8000 1.1350 0.9000 ;
      RECT 0.2400 0.9900 0.3300 1.4700 ;
      RECT 0.8150 0.5300 0.9050 0.9000 ;
      RECT 0.5850 1.5600 0.7650 1.9600 ;
      RECT 0.2400 1.4700 0.7650 1.5600 ;
      RECT 0.6750 0.9900 0.7650 1.4700 ;
      RECT 1.4850 1.3550 1.5750 1.5850 ;
      RECT 1.2350 1.2650 1.5750 1.3550 ;
      RECT 1.2350 1.2050 1.3250 1.2650 ;
      RECT 0.8550 1.1150 1.3250 1.2050 ;
      RECT 1.2350 0.6350 1.3250 1.1150 ;
      RECT 1.2350 0.5450 1.6450 0.6350 ;
      RECT 1.9450 0.6600 2.0350 1.7200 ;
      RECT 2.1250 1.5000 2.7500 1.5900 ;
      RECT 2.6500 0.7100 2.7500 1.5000 ;
      RECT 2.5500 0.6200 2.7500 0.7100 ;
      RECT 1.4450 0.7450 1.5350 1.0850 ;
      RECT 1.7550 1.1750 1.8450 1.8300 ;
      RECT 1.4450 1.0850 1.8450 1.1750 ;
      RECT 1.7550 1.8300 2.2150 1.9200 ;
      RECT 2.1250 1.5900 2.2150 1.8300 ;
  END
END LATSQN_X1M_A12TH

MACRO LATSQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.5400 0.3200 0.6300 0.5450 ;
        RECT 1.0950 0.3200 1.1850 0.4650 ;
        RECT 2.5350 0.3200 2.6250 0.6250 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0350 0.5500 1.4800 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3050 1.2500 2.7300 1.3500 ;
    END
    ANTENNAGATEAREA 0.0558 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3550 0.8100 2.7500 0.9100 ;
        RECT 2.3550 0.5700 2.4450 0.8100 ;
        RECT 2.6500 0.9100 2.7500 1.0800 ;
        RECT 1.9150 0.4800 2.4450 0.5700 ;
        RECT 1.9150 0.5700 2.0050 1.0350 ;
        RECT 1.7850 1.0350 2.0050 1.1250 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9450 1.1500 1.3000 ;
        RECT 0.8750 1.3000 1.1500 1.4000 ;
        RECT 0.7800 0.8450 1.1500 0.9450 ;
        RECT 0.8750 1.4000 0.9650 1.6900 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.0800 1.7800 0.1700 2.0800 ;
        RECT 0.6150 1.7800 0.7050 2.0800 ;
        RECT 1.1350 1.7800 1.2250 2.0800 ;
        RECT 2.4950 1.7050 2.5850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0450 1.5900 0.7700 1.6800 ;
      RECT 0.6800 1.0700 0.7700 1.5900 ;
      RECT 0.3400 1.6800 0.4300 1.9750 ;
      RECT 0.0450 0.7800 0.1350 1.5900 ;
      RECT 0.0450 0.4100 0.1700 0.7800 ;
      RECT 1.7300 1.5350 1.8200 1.9200 ;
      RECT 1.3850 1.4450 1.8200 1.5350 ;
      RECT 0.4550 0.6350 1.8200 0.7250 ;
      RECT 1.7300 0.5150 1.8200 0.6350 ;
      RECT 1.3850 0.7250 1.4750 1.4450 ;
      RECT 0.4550 0.7250 0.5450 0.8300 ;
      RECT 0.2450 0.8300 0.5450 0.9200 ;
      RECT 0.2450 0.9200 0.3350 1.5000 ;
      RECT 2.0950 0.7700 2.1850 1.7200 ;
      RECT 2.0950 0.6800 2.2650 0.7700 ;
      RECT 2.2950 1.5050 2.9400 1.5950 ;
      RECT 2.8300 1.5950 2.9400 1.9050 ;
      RECT 2.8500 0.7050 2.9400 1.5050 ;
      RECT 2.8300 0.4950 2.9400 0.7050 ;
      RECT 1.5650 0.8350 1.6550 1.2450 ;
      RECT 1.9100 1.3350 2.0000 1.8300 ;
      RECT 1.5650 1.2450 2.0000 1.3350 ;
      RECT 1.9100 1.8300 2.3850 1.9200 ;
      RECT 2.2950 1.5950 2.3850 1.8300 ;
  END
END LATSQN_X2M_A12TH

MACRO LATSQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6650 ;
        RECT 0.8600 0.3200 0.9500 0.6650 ;
        RECT 1.5800 0.3200 1.6700 0.5800 ;
        RECT 2.7700 0.3200 2.8600 0.8250 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0150 1.1050 1.1500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5950 1.1900 2.7500 1.4000 ;
        RECT 2.6500 1.4000 2.7500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0250 2.9500 1.1900 ;
        RECT 2.5900 0.9350 2.9500 1.0250 ;
        RECT 2.5900 0.5700 2.6800 0.9350 ;
        RECT 2.2300 0.4800 2.6800 0.5700 ;
        RECT 2.2300 0.5700 2.3200 0.9250 ;
        RECT 2.1900 0.9250 2.3200 1.0950 ;
    END
    ANTENNAGATEAREA 0.0816 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4500 0.6900 1.5500 ;
        RECT 0.0800 1.5500 0.1700 1.8400 ;
        RECT 0.6000 1.5500 0.6900 1.8400 ;
        RECT 0.0800 0.9500 0.1800 1.4500 ;
        RECT 0.0800 0.8500 0.6900 0.9500 ;
        RECT 0.0800 0.5600 0.1700 0.8500 ;
        RECT 0.6000 0.5600 0.6900 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.7000 2.0100 2.7900 2.0800 ;
        RECT 0.3400 1.8200 0.4300 2.0800 ;
        RECT 0.8600 1.8200 0.9500 2.0800 ;
        RECT 1.3800 1.8200 1.4700 2.0800 ;
        RECT 1.5800 1.5650 1.6700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.2400 1.0450 1.6250 1.1450 ;
      RECT 1.1200 1.6250 1.2100 1.9450 ;
      RECT 1.1200 1.6200 1.3300 1.6250 ;
      RECT 0.7900 1.5300 1.3300 1.6200 ;
      RECT 1.2400 1.1450 1.3300 1.5300 ;
      RECT 0.7900 1.1800 0.8800 1.5300 ;
      RECT 0.3050 1.0900 0.8800 1.1800 ;
      RECT 1.3500 0.5600 1.4400 1.0450 ;
      RECT 2.0500 1.4750 2.1400 1.7550 ;
      RECT 1.4200 1.3850 2.1400 1.4750 ;
      RECT 1.7150 0.7600 1.8050 1.3850 ;
      RECT 1.7150 0.6700 2.1200 0.7600 ;
      RECT 2.0300 0.4100 2.1200 0.6700 ;
      RECT 1.4200 1.2700 1.5100 1.3850 ;
      RECT 2.4100 0.6800 2.5000 1.7200 ;
      RECT 3.0300 1.9200 3.1300 1.9700 ;
      RECT 2.2300 1.8300 3.1300 1.9200 ;
      RECT 3.0300 1.5600 3.1300 1.8300 ;
      RECT 3.0400 0.8600 3.1300 1.5600 ;
      RECT 3.0300 0.4500 3.1300 0.8600 ;
      RECT 1.9250 0.8500 2.0150 1.2050 ;
      RECT 2.2300 1.2950 2.3200 1.8300 ;
      RECT 1.9250 1.2050 2.3200 1.2950 ;
  END
END LATSQN_X3M_A12TH

MACRO LATSQN_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3450 0.3200 0.4950 0.3800 ;
        RECT 1.6800 0.3200 1.7700 0.6300 ;
        RECT 2.6150 0.3200 2.7050 0.6300 ;
        RECT 3.1700 0.3200 3.2600 0.6650 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0500 0.5550 1.5300 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6100 1.0500 2.6250 1.1500 ;
    END
    ANTENNAGATEAREA 0.162 ;
  END SN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9100 1.4500 3.5200 1.5500 ;
        RECT 2.9100 1.5500 3.0000 1.8600 ;
        RECT 3.4300 1.5500 3.5200 1.8600 ;
        RECT 3.4200 0.9500 3.5200 1.4500 ;
        RECT 2.9100 0.8500 3.5200 0.9500 ;
        RECT 2.9100 0.5600 3.0000 0.8500 ;
        RECT 3.4300 0.5600 3.5200 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.3150 2.0550 0.5250 2.0800 ;
        RECT 1.6100 1.7700 1.7000 2.0800 ;
        RECT 2.1300 1.7700 2.2200 2.0800 ;
        RECT 2.6500 1.7700 2.7400 2.0800 ;
        RECT 3.1700 1.7700 3.2600 2.0800 ;
    END
  END VDD

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.5700 0.9500 1.2000 ;
        RECT 0.4500 0.4800 0.9500 0.5700 ;
        RECT 0.4500 0.5700 0.5500 0.8500 ;
        RECT 0.2350 0.8500 0.5500 0.9400 ;
        RECT 0.2350 0.9400 0.3250 1.1200 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END G
  OBS
    LAYER M1 ;
      RECT 0.6450 0.6800 0.7350 1.6900 ;
      RECT 0.0550 1.8300 0.9450 1.9200 ;
      RECT 0.8550 1.4200 0.9450 1.8300 ;
      RECT 0.8550 1.3300 1.1750 1.4200 ;
      RECT 1.0850 1.0950 1.1750 1.3300 ;
      RECT 1.0850 1.0050 1.2650 1.0950 ;
      RECT 1.1750 0.7550 1.2650 1.0050 ;
      RECT 0.0550 1.7100 0.1700 1.8300 ;
      RECT 0.0550 0.7800 0.1450 1.7100 ;
      RECT 0.0550 0.4100 0.1700 0.7800 ;
      RECT 1.2650 1.2400 2.3800 1.3300 ;
      RECT 1.0400 1.6200 1.1300 1.9600 ;
      RECT 1.0400 1.5300 1.3550 1.6200 ;
      RECT 1.2650 1.3300 1.3550 1.5300 ;
      RECT 1.3900 0.6450 1.4800 1.2400 ;
      RECT 1.0400 0.5550 1.4800 0.6450 ;
      RECT 1.0400 0.4300 1.1300 0.5550 ;
      RECT 2.7300 1.0900 3.1650 1.1800 ;
      RECT 1.4650 1.4200 2.8200 1.5100 ;
      RECT 2.7300 1.1800 2.8200 1.4200 ;
      RECT 2.7300 0.9300 2.8200 1.0900 ;
      RECT 2.1300 0.8400 2.8200 0.9300 ;
      RECT 1.8700 1.5100 1.9600 1.9700 ;
      RECT 2.3900 1.5100 2.4800 1.9700 ;
      RECT 2.1300 0.5200 2.2200 0.8400 ;
  END
END LATSQN_X4M_A12TH

MACRO M2DFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4250 0.3200 0.5250 0.8050 ;
        RECT 1.5800 0.3200 1.7500 0.3750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8200 0.9100 5.9700 1.3000 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.7550 5.1500 1.3150 ;
        RECT 5.0500 1.3150 5.1900 1.7200 ;
        RECT 5.0500 0.6650 5.2300 0.7550 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8650 1.5700 1.2550 ;
    END
    ANTENNAGATEAREA 0.0324 ;
  END D0

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8550 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END S0

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.8500 0.7500 1.2650 ;
    END
    ANTENNAGATEAREA 0.0324 ;
  END D1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.6300 2.0200 5.8000 2.0800 ;
        RECT 0.4000 1.7500 0.5100 2.0800 ;
        RECT 1.6300 1.4500 1.7300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7050 1.3800 0.9400 1.4700 ;
      RECT 0.8400 0.7400 0.9400 1.3800 ;
      RECT 0.6750 0.6500 0.9400 0.7400 ;
      RECT 0.6800 1.6500 1.1050 1.7350 ;
      RECT 0.0500 1.6450 1.1050 1.6500 ;
      RECT 0.0500 1.5600 0.7700 1.6450 ;
      RECT 0.0500 1.4350 0.1700 1.5600 ;
      RECT 0.0500 0.7550 0.1400 1.4350 ;
      RECT 0.0500 0.6650 0.2400 0.7550 ;
      RECT 1.3750 1.4450 1.4650 1.6100 ;
      RECT 1.2300 1.3550 1.4650 1.4450 ;
      RECT 1.2300 0.7600 1.3200 1.3550 ;
      RECT 1.2300 0.6700 1.4400 0.7600 ;
      RECT 1.0300 0.4900 1.8600 0.5800 ;
      RECT 1.7700 0.5800 1.8600 1.2750 ;
      RECT 1.0300 0.5800 1.1200 1.5350 ;
      RECT 1.9500 0.6050 2.0400 1.6400 ;
      RECT 2.1750 1.5000 2.4200 1.5900 ;
      RECT 2.3300 0.7700 2.4200 1.5000 ;
      RECT 2.3300 0.6800 3.1250 0.7700 ;
      RECT 3.0350 0.7700 3.1250 1.3000 ;
      RECT 2.6250 1.4750 3.3250 1.5650 ;
      RECT 2.6250 1.1650 2.7150 1.4750 ;
      RECT 3.2350 0.7700 3.3250 1.4750 ;
      RECT 3.2350 0.6800 3.4100 0.7700 ;
      RECT 3.4300 1.4800 3.9750 1.5700 ;
      RECT 3.8850 0.7700 3.9750 1.4800 ;
      RECT 3.6800 0.6800 4.4400 0.7700 ;
      RECT 4.3500 0.7700 4.4400 1.2950 ;
      RECT 4.0850 1.4900 4.8200 1.5800 ;
      RECT 4.7300 1.1750 4.8200 1.4900 ;
      RECT 4.0850 0.9700 4.1750 1.4900 ;
      RECT 4.7300 1.0850 4.9500 1.1750 ;
      RECT 4.7300 0.7700 4.8200 1.0850 ;
      RECT 4.5500 0.6800 4.8200 0.7700 ;
      RECT 2.1500 0.4800 5.4400 0.5700 ;
      RECT 5.3500 0.5700 5.4400 1.6300 ;
      RECT 3.5000 1.2800 3.7650 1.3700 ;
      RECT 3.5000 0.5700 3.5900 1.2800 ;
      RECT 2.1500 0.5700 2.2400 1.3850 ;
      RECT 2.4250 0.4100 2.5950 0.4800 ;
      RECT 5.5300 1.5000 6.1350 1.5900 ;
      RECT 5.5300 0.6400 6.1350 0.7300 ;
      RECT 2.2850 1.8300 5.6200 1.9200 ;
      RECT 5.5300 1.5900 5.6200 1.8300 ;
      RECT 5.5300 0.7300 5.6200 1.5000 ;
  END
END M2DFFQN_X0P5M_A12TH

MACRO M2DFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4050 0.3200 0.5050 0.7150 ;
        RECT 1.5800 0.3200 1.7500 0.3750 ;
    END
  END VSS

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8650 1.5700 1.2550 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END D0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.6300 2.0200 5.8000 2.0800 ;
        RECT 0.3700 1.7500 0.5400 2.0800 ;
        RECT 1.6300 1.4050 1.7300 2.0800 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.7550 5.1500 1.3150 ;
        RECT 5.0500 1.3150 5.1950 1.4150 ;
        RECT 5.0500 0.6650 5.2300 0.7550 ;
        RECT 5.0950 1.4150 5.1950 1.7200 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8200 0.9100 5.9700 1.3000 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CK

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0702 ;
  END S0

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 0.7050 1.3800 0.9400 1.4700 ;
      RECT 0.8400 0.6750 0.9400 1.3800 ;
      RECT 0.7050 0.5850 0.9400 0.6750 ;
      RECT 0.7850 1.6950 1.1050 1.7850 ;
      RECT 0.7850 1.6500 0.8750 1.6950 ;
      RECT 0.0500 1.5600 0.8750 1.6500 ;
      RECT 0.0500 1.4400 0.1700 1.5600 ;
      RECT 0.0500 0.6950 0.1400 1.4400 ;
      RECT 0.0500 0.5750 0.2350 0.6950 ;
      RECT 1.3750 1.4600 1.4650 1.7850 ;
      RECT 1.2250 1.3700 1.4650 1.4600 ;
      RECT 1.2250 0.7600 1.3150 1.3700 ;
      RECT 1.2250 0.6700 1.4400 0.7600 ;
      RECT 1.0300 0.4900 1.8600 0.5800 ;
      RECT 1.7700 0.5800 1.8600 1.2750 ;
      RECT 1.0300 0.5800 1.1200 1.5750 ;
      RECT 1.9500 0.5650 2.0400 1.6650 ;
      RECT 2.1750 1.5000 2.4200 1.5900 ;
      RECT 2.3300 0.7700 2.4200 1.5000 ;
      RECT 2.3300 0.6800 3.1250 0.7700 ;
      RECT 3.0350 0.7700 3.1250 1.2750 ;
      RECT 2.6250 1.4800 3.3250 1.5700 ;
      RECT 2.6250 1.1650 2.7150 1.4800 ;
      RECT 3.2350 0.7700 3.3250 1.4800 ;
      RECT 3.2350 0.6800 3.4100 0.7700 ;
      RECT 3.4800 1.5900 3.9750 1.6800 ;
      RECT 3.8850 0.7700 3.9750 1.5900 ;
      RECT 3.6800 0.6800 4.4400 0.7700 ;
      RECT 4.3500 0.7700 4.4400 0.9700 ;
      RECT 4.3500 0.9700 4.5300 1.0600 ;
      RECT 4.4400 1.0600 4.5300 1.4000 ;
      RECT 4.0850 1.6350 4.7250 1.7250 ;
      RECT 4.6350 1.1550 4.7250 1.6350 ;
      RECT 4.0850 1.0500 4.1750 1.6350 ;
      RECT 4.6350 1.0650 4.9400 1.1550 ;
      RECT 4.6350 0.7550 4.7250 1.0650 ;
      RECT 4.5500 0.6650 4.7250 0.7550 ;
      RECT 2.1500 0.4800 5.4400 0.5700 ;
      RECT 5.3500 0.5700 5.4400 1.6100 ;
      RECT 3.6750 1.0350 3.7650 1.4550 ;
      RECT 3.5000 0.9450 3.7650 1.0350 ;
      RECT 3.5000 0.5700 3.5900 0.9450 ;
      RECT 2.1500 0.5700 2.2400 1.3850 ;
      RECT 2.4250 0.4100 2.5950 0.4800 ;
      RECT 5.5300 1.4800 6.1150 1.5700 ;
      RECT 5.5300 0.6300 6.1150 0.7200 ;
      RECT 2.2850 1.8300 5.6200 1.9200 ;
      RECT 5.5300 1.5700 5.6200 1.8300 ;
      RECT 5.5300 0.7200 5.6200 1.4800 ;
  END
END M2DFFQN_X1M_A12TH

MACRO M2DFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7200 ;
        RECT 2.7450 0.3200 2.9150 0.3800 ;
        RECT 5.7300 0.3200 5.9000 0.5050 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9050 0.5500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END S0

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.8350 5.9550 1.2600 ;
    END
    ANTENNAGATEAREA 0.033 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8100 5.1500 1.2550 ;
        RECT 4.9100 1.2550 5.1500 1.3550 ;
        RECT 4.8500 0.7100 5.1500 0.8100 ;
        RECT 4.9100 1.3550 5.0100 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 3.9050 2.0200 4.2750 2.0800 ;
        RECT 2.5750 2.0150 2.9450 2.0800 ;
        RECT 0.3150 1.8700 0.4850 2.0800 ;
        RECT 1.5800 1.4600 1.6800 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 0.8650 1.5500 1.2750 ;
    END
    ANTENNAGATEAREA 0.0462 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 0.6400 0.7250 0.7300 1.5800 ;
      RECT 0.6000 0.5550 0.7300 0.7250 ;
      RECT 0.0550 1.6900 0.9100 1.7800 ;
      RECT 0.8200 1.1400 0.9100 1.6900 ;
      RECT 0.2550 0.9000 0.3450 1.6900 ;
      RECT 0.0950 0.8100 0.3450 0.9000 ;
      RECT 0.0950 0.4300 0.1850 0.8100 ;
      RECT 1.2600 0.7550 1.3500 1.7750 ;
      RECT 1.1550 0.6650 1.3500 0.7550 ;
      RECT 0.8900 0.4800 1.8150 0.5700 ;
      RECT 1.7250 0.5700 1.8150 1.3150 ;
      RECT 1.0000 0.9150 1.0900 1.7750 ;
      RECT 0.8900 0.8250 1.0900 0.9150 ;
      RECT 0.8900 0.5700 0.9800 0.8250 ;
      RECT 1.9050 0.4450 1.9950 1.8050 ;
      RECT 2.1400 1.5250 2.3950 1.6150 ;
      RECT 2.3050 0.7500 2.3950 1.5250 ;
      RECT 2.3050 0.6600 3.0100 0.7500 ;
      RECT 2.9200 0.7500 3.0100 1.3300 ;
      RECT 2.6100 1.5700 3.2100 1.6600 ;
      RECT 2.6100 1.0250 2.7000 1.5700 ;
      RECT 3.1200 0.6600 3.2100 1.5700 ;
      RECT 3.4800 1.6300 3.9150 1.7200 ;
      RECT 3.8250 0.7500 3.9150 1.6300 ;
      RECT 3.5150 0.6600 4.2750 0.7500 ;
      RECT 3.5150 0.7500 3.6150 0.8600 ;
      RECT 4.1850 0.7500 4.2750 1.0900 ;
      RECT 4.1850 1.0900 4.3750 1.1800 ;
      RECT 4.4000 1.3900 4.5000 1.7150 ;
      RECT 4.0050 1.3000 4.6750 1.3900 ;
      RECT 4.5850 1.1650 4.6750 1.3000 ;
      RECT 4.0050 1.0400 4.0950 1.3000 ;
      RECT 4.5850 1.0650 4.8450 1.1650 ;
      RECT 4.5850 0.9350 4.6750 1.0650 ;
      RECT 4.3650 0.8350 4.6750 0.9350 ;
      RECT 2.1250 0.4800 5.5150 0.5700 ;
      RECT 5.4250 0.5700 5.5150 1.6500 ;
      RECT 3.6250 1.0700 3.7150 1.5050 ;
      RECT 3.3300 0.9800 3.7150 1.0700 ;
      RECT 3.3300 0.5700 3.4200 0.9800 ;
      RECT 2.1250 0.5700 2.2150 1.4050 ;
      RECT 2.3700 0.4250 2.5400 0.4800 ;
      RECT 2.3700 1.8300 6.1200 1.9200 ;
      RECT 6.0300 1.4900 6.1200 1.8300 ;
      RECT 5.6150 0.6100 6.1200 0.7000 ;
      RECT 6.0300 0.4450 6.1200 0.6100 ;
      RECT 5.6150 0.7000 5.7050 1.8300 ;
      RECT 3.3000 1.3750 3.3900 1.8300 ;
      RECT 3.3000 1.2050 3.4400 1.3750 ;
  END
END M2DFFQN_X2M_A12TH

MACRO M2DFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.7200 ;
        RECT 2.7450 0.3200 2.9150 0.3800 ;
        RECT 5.9300 0.3200 6.1000 0.5050 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9050 0.5500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END S0

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.8350 6.1550 1.2600 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8800 1.2500 5.5000 1.3500 ;
        RECT 4.8800 1.3500 4.9800 1.7200 ;
        RECT 5.4000 1.3500 5.5000 1.7250 ;
        RECT 5.4000 0.8100 5.5000 1.2500 ;
        RECT 4.8200 0.7100 5.5000 0.8100 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 2.5750 2.0250 2.9450 2.0800 ;
        RECT 0.3150 1.8700 0.4850 2.0800 ;
        RECT 1.5800 1.5300 1.6800 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 0.8600 1.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 0.6400 0.7250 0.7300 1.5800 ;
      RECT 0.6000 0.5550 0.7300 0.7250 ;
      RECT 0.0550 1.6900 0.9100 1.7800 ;
      RECT 0.8200 1.1400 0.9100 1.6900 ;
      RECT 0.2550 0.9000 0.3450 1.6900 ;
      RECT 0.0950 0.8100 0.3450 0.9000 ;
      RECT 0.0950 0.4400 0.1850 0.8100 ;
      RECT 1.2600 0.7550 1.3500 1.8150 ;
      RECT 1.1550 0.6650 1.3500 0.7550 ;
      RECT 0.8900 0.4800 1.8250 0.5700 ;
      RECT 1.7350 0.5700 1.8250 1.3150 ;
      RECT 1.0000 0.9150 1.0900 1.8150 ;
      RECT 0.8900 0.8250 1.0900 0.9150 ;
      RECT 0.8900 0.5700 0.9800 0.8250 ;
      RECT 1.9400 0.4450 2.0300 1.8850 ;
      RECT 2.1400 1.5250 2.3950 1.6150 ;
      RECT 2.3050 0.7500 2.3950 1.5250 ;
      RECT 2.3050 0.6600 3.0100 0.7500 ;
      RECT 2.9200 0.7500 3.0100 1.3300 ;
      RECT 2.6100 1.6150 3.2100 1.7050 ;
      RECT 2.6100 1.0250 2.7000 1.6150 ;
      RECT 3.1200 0.6600 3.2100 1.6150 ;
      RECT 3.4800 1.6300 3.8850 1.7200 ;
      RECT 3.7950 0.7500 3.8850 1.6300 ;
      RECT 3.5150 0.6600 4.2450 0.7500 ;
      RECT 3.5150 0.7500 3.6150 0.8600 ;
      RECT 4.1550 0.7500 4.2450 1.0900 ;
      RECT 4.1550 1.0900 4.3450 1.1800 ;
      RECT 4.4350 1.0700 5.1700 1.1600 ;
      RECT 4.3700 1.3900 4.4700 1.7150 ;
      RECT 3.9750 1.3000 4.5250 1.3900 ;
      RECT 4.4350 1.1600 4.5250 1.3000 ;
      RECT 3.9750 1.0400 4.0650 1.3000 ;
      RECT 4.4350 0.9300 4.5250 1.0700 ;
      RECT 4.3350 0.8400 4.5250 0.9300 ;
      RECT 2.1250 0.4800 5.7450 0.5700 ;
      RECT 5.6550 0.5700 5.7450 1.7200 ;
      RECT 3.6150 1.0700 3.7050 1.5200 ;
      RECT 3.3300 0.9800 3.7050 1.0700 ;
      RECT 3.3300 0.5700 3.4200 0.9800 ;
      RECT 2.1250 0.5700 2.2150 1.4050 ;
      RECT 2.3700 0.4250 2.5400 0.4800 ;
      RECT 2.3700 1.8300 6.3200 1.9200 ;
      RECT 6.2300 1.3400 6.3200 1.8300 ;
      RECT 5.8350 0.6100 6.3200 0.7000 ;
      RECT 6.2300 0.4450 6.3200 0.6100 ;
      RECT 5.8350 0.7000 5.9250 1.8300 ;
      RECT 3.3000 1.3750 3.3900 1.8300 ;
      RECT 3.3000 1.2050 3.4400 1.3750 ;
  END
END M2DFFQN_X3M_A12TH

MACRO M2DFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4250 0.3200 0.5250 0.7400 ;
        RECT 1.5800 0.3200 1.7500 0.3750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8200 0.9100 5.9500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8150 5.1500 1.3150 ;
        RECT 5.0500 1.3150 5.1950 1.4150 ;
        RECT 5.0500 0.7150 5.2500 0.8150 ;
        RECT 5.0950 1.4150 5.1950 1.7200 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8650 1.5700 1.2550 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END D0

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8100 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END S0

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.8100 0.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END D1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.6300 2.0200 5.8000 2.0800 ;
        RECT 0.3700 1.7500 0.5400 2.0800 ;
        RECT 1.6300 1.4650 1.7300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7050 1.3800 0.9400 1.4700 ;
      RECT 0.8400 0.7000 0.9400 1.3800 ;
      RECT 0.6750 0.6100 0.9400 0.7000 ;
      RECT 0.7850 1.8800 1.1200 1.9700 ;
      RECT 0.7850 1.6500 0.8750 1.8800 ;
      RECT 0.0500 1.5600 0.8750 1.6500 ;
      RECT 0.0500 1.4650 0.1700 1.5600 ;
      RECT 0.0500 0.7150 0.1400 1.4650 ;
      RECT 0.0500 0.6250 0.2400 0.7150 ;
      RECT 1.3750 1.5900 1.4650 1.6750 ;
      RECT 1.2250 1.5000 1.4650 1.5900 ;
      RECT 1.2250 0.7600 1.3150 1.5000 ;
      RECT 1.2250 0.6700 1.4400 0.7600 ;
      RECT 1.0300 0.4900 1.8600 0.5800 ;
      RECT 1.7700 0.5800 1.8600 1.2900 ;
      RECT 1.0300 0.5800 1.1200 1.5450 ;
      RECT 1.9500 0.6050 2.0400 1.6400 ;
      RECT 2.1750 1.5000 2.4200 1.5900 ;
      RECT 2.3300 0.7700 2.4200 1.5000 ;
      RECT 2.3300 0.6800 3.1250 0.7700 ;
      RECT 3.0350 0.7700 3.1250 1.2950 ;
      RECT 2.6250 1.4750 3.3250 1.5650 ;
      RECT 2.6250 1.1650 2.7150 1.4750 ;
      RECT 3.2350 0.7700 3.3250 1.4750 ;
      RECT 3.2350 0.6800 3.4100 0.7700 ;
      RECT 4.5950 1.5650 4.6850 1.6250 ;
      RECT 4.0850 1.4750 4.6850 1.5650 ;
      RECT 4.0850 0.9700 4.1750 1.4750 ;
      RECT 4.5950 0.9500 4.6850 1.4750 ;
      RECT 4.5500 0.8600 4.7450 0.9500 ;
      RECT 3.4150 1.4800 3.9750 1.5700 ;
      RECT 3.8850 0.7700 3.9750 1.4800 ;
      RECT 3.6800 0.6800 4.9450 0.7700 ;
      RECT 4.3500 0.7700 4.4400 1.2950 ;
      RECT 4.8550 0.7700 4.9450 1.1500 ;
      RECT 2.1500 0.4800 5.4400 0.5700 ;
      RECT 5.3500 0.5700 5.4400 1.6300 ;
      RECT 3.5000 1.2800 3.7650 1.3700 ;
      RECT 3.5000 0.5700 3.5900 1.2800 ;
      RECT 2.1500 0.5700 2.2400 1.3900 ;
      RECT 2.4250 0.4100 2.5950 0.4800 ;
      RECT 5.5300 1.5000 6.1350 1.5900 ;
      RECT 5.5300 0.6400 6.1350 0.7300 ;
      RECT 2.2850 1.8300 5.6200 1.9200 ;
      RECT 5.5300 1.5900 5.6200 1.8300 ;
      RECT 5.5300 0.7300 5.6200 1.5000 ;
  END
END M2DFFQ_X0P5M_A12TH

MACRO M2DFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4050 0.3200 0.5050 0.7150 ;
        RECT 1.5800 0.3200 1.7500 0.3750 ;
    END
  END VSS

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8500 1.5700 1.2550 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END D0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.6500 2.0200 5.8200 2.0800 ;
        RECT 0.3700 1.8500 0.5400 2.0800 ;
        RECT 1.6300 1.4550 1.7300 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.7800 5.1500 1.3150 ;
        RECT 5.0500 1.3150 5.1950 1.4150 ;
        RECT 5.0500 0.6800 5.2500 0.7800 ;
        RECT 5.0950 1.4150 5.1950 1.7200 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8300 0.9100 5.9500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END CK

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END S0

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 0.7050 1.3800 0.9400 1.4700 ;
      RECT 0.8400 0.6750 0.9400 1.3800 ;
      RECT 0.7050 0.5850 0.9400 0.6750 ;
      RECT 0.7850 1.8800 1.1200 1.9700 ;
      RECT 0.7850 1.7400 0.8750 1.8800 ;
      RECT 0.0500 1.6500 0.8750 1.7400 ;
      RECT 0.0800 1.7400 0.1700 1.8400 ;
      RECT 0.0500 0.6950 0.1400 1.6500 ;
      RECT 0.0500 0.5750 0.2350 0.6950 ;
      RECT 1.3750 1.5600 1.4650 1.8400 ;
      RECT 1.2100 1.4700 1.4650 1.5600 ;
      RECT 1.2100 0.7600 1.3000 1.4700 ;
      RECT 1.2100 0.6700 1.4400 0.7600 ;
      RECT 1.0300 0.4900 1.8600 0.5800 ;
      RECT 1.7700 0.5800 1.8600 1.2750 ;
      RECT 1.0300 0.5800 1.1200 1.5750 ;
      RECT 1.9500 0.5650 2.0400 1.6650 ;
      RECT 2.1750 1.5000 2.4200 1.5900 ;
      RECT 2.3300 0.7700 2.4200 1.5000 ;
      RECT 2.3300 0.6800 3.1250 0.7700 ;
      RECT 3.0350 0.7700 3.1250 1.2950 ;
      RECT 2.6250 1.4750 3.3250 1.5650 ;
      RECT 2.6250 1.1650 2.7150 1.4750 ;
      RECT 3.2350 0.7700 3.3250 1.4750 ;
      RECT 3.2350 0.6800 3.4100 0.7700 ;
      RECT 4.0850 1.6350 4.7250 1.7250 ;
      RECT 4.0850 1.0850 4.1750 1.6350 ;
      RECT 4.6350 0.9500 4.7250 1.6350 ;
      RECT 4.5500 0.8600 4.7250 0.9500 ;
      RECT 3.4100 1.6400 3.9750 1.7300 ;
      RECT 3.8850 0.7700 3.9750 1.6400 ;
      RECT 3.6800 0.6800 4.9200 0.7700 ;
      RECT 4.3500 0.7700 4.4400 1.2950 ;
      RECT 4.8300 0.7700 4.9200 1.1500 ;
      RECT 2.1500 0.4800 5.4500 0.5700 ;
      RECT 5.3600 0.5700 5.4500 1.6100 ;
      RECT 3.6750 1.0350 3.7650 1.5300 ;
      RECT 3.5000 0.9450 3.7650 1.0350 ;
      RECT 3.5000 0.5700 3.5900 0.9450 ;
      RECT 2.1500 0.5700 2.2400 1.3900 ;
      RECT 2.4250 0.4100 2.5950 0.4800 ;
      RECT 5.5400 1.5000 6.1350 1.5900 ;
      RECT 5.5400 0.6300 6.1350 0.7200 ;
      RECT 2.2850 1.8300 5.6400 1.9200 ;
      RECT 5.5400 1.5900 5.6300 1.8300 ;
      RECT 5.5400 0.7200 5.6300 1.5000 ;
      RECT 3.3550 1.9200 3.5250 1.9650 ;
  END
END M2DFFQ_X1M_A12TH

MACRO M2DFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6900 ;
        RECT 1.5000 0.3200 1.6700 0.3900 ;
        RECT 2.7950 0.3200 2.9650 0.3300 ;
        RECT 5.7300 0.3200 5.9000 0.5050 ;
    END
  END VSS

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0474 ;
  END D0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.3150 1.8800 0.4850 2.0800 ;
        RECT 1.6600 1.5000 1.7500 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8850 5.1500 1.2500 ;
        RECT 4.9150 1.2500 5.1500 1.3500 ;
        RECT 4.8600 0.7850 5.1500 0.8850 ;
        RECT 4.9150 1.3500 5.0050 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.8350 5.9500 1.2600 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END CK

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END S0

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0474 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 0.6400 0.6900 0.7300 1.6000 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0550 1.7000 0.9300 1.7900 ;
      RECT 0.8400 1.0600 0.9300 1.7000 ;
      RECT 0.2550 0.8700 0.3450 1.7000 ;
      RECT 0.0950 0.7800 0.3450 0.8700 ;
      RECT 0.0950 0.4800 0.1850 0.7800 ;
      RECT 1.2700 1.4600 1.3700 1.6850 ;
      RECT 1.2700 0.7550 1.3600 1.4600 ;
      RECT 1.0950 0.6650 1.3600 0.7550 ;
      RECT 0.8900 0.4800 1.8450 0.5700 ;
      RECT 1.7550 0.5700 1.8450 1.1000 ;
      RECT 1.0200 0.9500 1.1100 1.6850 ;
      RECT 0.8900 0.8600 1.1100 0.9500 ;
      RECT 0.8900 0.5700 0.9800 0.8600 ;
      RECT 1.9400 0.4800 2.0300 1.9000 ;
      RECT 2.2000 1.6000 2.2900 1.9350 ;
      RECT 2.2000 1.5100 2.3950 1.6000 ;
      RECT 2.3050 0.7550 2.3950 1.5100 ;
      RECT 2.3050 0.6650 3.0100 0.7550 ;
      RECT 2.9200 0.7550 3.0100 1.1750 ;
      RECT 2.6100 1.5700 3.2100 1.6600 ;
      RECT 2.6100 1.1150 2.7000 1.5700 ;
      RECT 3.1200 0.6600 3.2100 1.5700 ;
      RECT 4.0050 1.5300 4.5550 1.6200 ;
      RECT 4.0050 1.0400 4.0950 1.5300 ;
      RECT 4.4650 0.9500 4.5550 1.5300 ;
      RECT 4.3650 0.8600 4.5550 0.9500 ;
      RECT 3.4800 1.5450 3.9150 1.6350 ;
      RECT 3.8250 0.7500 3.9150 1.5450 ;
      RECT 3.5200 0.6600 4.7650 0.7500 ;
      RECT 3.5200 0.7500 3.6100 0.8350 ;
      RECT 4.1850 0.7500 4.2750 1.1050 ;
      RECT 4.6750 0.7500 4.7650 1.2200 ;
      RECT 4.1850 1.1050 4.3750 1.1950 ;
      RECT 5.4050 1.3500 5.5300 1.5300 ;
      RECT 5.4400 0.6650 5.5300 1.3500 ;
      RECT 5.4250 0.5700 5.5300 0.6650 ;
      RECT 2.1250 0.4800 5.5300 0.5700 ;
      RECT 2.1250 0.5700 2.2150 1.4000 ;
      RECT 3.3300 0.5700 3.4200 0.9550 ;
      RECT 2.3700 0.4250 2.5400 0.4800 ;
      RECT 3.3300 0.9550 3.7050 1.0450 ;
      RECT 3.6150 1.0450 3.7050 1.4550 ;
      RECT 5.4100 1.6450 6.1200 1.7350 ;
      RECT 6.0300 1.5000 6.1200 1.6450 ;
      RECT 5.6200 0.6100 6.1200 0.7000 ;
      RECT 6.0300 0.4450 6.1200 0.6100 ;
      RECT 2.3800 1.8300 5.5000 1.9200 ;
      RECT 5.4100 1.7350 5.5000 1.8300 ;
      RECT 5.6200 0.7000 5.7100 1.6450 ;
      RECT 3.3000 1.3850 3.3900 1.8300 ;
      RECT 3.3000 1.2150 3.4400 1.3850 ;
  END
END M2DFFQ_X2M_A12TH

MACRO M2DFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6900 ;
        RECT 5.9300 0.3200 6.1000 0.5050 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END S0

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.8350 6.1550 1.2600 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8350 1.0500 5.4550 1.1500 ;
        RECT 4.8350 1.1500 4.9350 1.7300 ;
        RECT 5.3550 1.1500 5.4550 1.7200 ;
        RECT 4.8350 0.7000 4.9350 1.0500 ;
        RECT 5.3650 0.7000 5.4550 1.0500 ;
    END
    ANTENNADIFFAREA 0.595725 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.3150 1.8800 0.4850 2.0800 ;
        RECT 1.6600 1.5000 1.7500 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8600 1.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D0
  OBS
    LAYER M1 ;
      RECT 0.6400 0.6900 0.7300 1.5800 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0550 1.7000 0.9100 1.7900 ;
      RECT 0.8200 1.1050 0.9100 1.7000 ;
      RECT 0.2550 0.8900 0.3450 1.7000 ;
      RECT 0.0950 0.8000 0.3450 0.8900 ;
      RECT 0.0950 0.4800 0.1850 0.8000 ;
      RECT 1.2600 1.1150 1.3500 1.6600 ;
      RECT 1.2100 1.0250 1.3500 1.1150 ;
      RECT 1.2100 0.7550 1.3000 1.0250 ;
      RECT 1.0950 0.6650 1.3000 0.7550 ;
      RECT 0.8900 0.4800 1.7950 0.5700 ;
      RECT 1.7050 0.5700 1.7950 1.1550 ;
      RECT 1.0000 0.9500 1.0900 1.6750 ;
      RECT 0.8900 0.8600 1.0900 0.9500 ;
      RECT 0.8900 0.5700 0.9800 0.8600 ;
      RECT 1.9400 0.4800 2.0300 1.8900 ;
      RECT 2.2000 1.5900 2.2900 1.9250 ;
      RECT 2.2000 1.5000 2.3950 1.5900 ;
      RECT 2.3050 0.7550 2.3950 1.5000 ;
      RECT 2.3050 0.6650 2.9650 0.7550 ;
      RECT 2.8750 0.7550 2.9650 1.1000 ;
      RECT 3.0550 1.3000 3.1450 1.6600 ;
      RECT 2.5500 1.2100 3.1450 1.3000 ;
      RECT 3.0550 0.8900 3.1450 1.2100 ;
      RECT 3.0550 0.6800 3.1800 0.8900 ;
      RECT 3.9300 1.5300 4.4800 1.6200 ;
      RECT 3.9300 1.0400 4.0200 1.5300 ;
      RECT 4.3900 0.9500 4.4800 1.5300 ;
      RECT 4.2900 0.8600 4.4800 0.9500 ;
      RECT 3.4150 1.5550 3.8400 1.6450 ;
      RECT 3.7500 0.7500 3.8400 1.5550 ;
      RECT 3.4550 0.6600 4.6900 0.7500 ;
      RECT 3.4550 0.7500 3.5450 0.8450 ;
      RECT 4.1100 0.7500 4.2000 1.1050 ;
      RECT 4.6000 0.7500 4.6900 1.2250 ;
      RECT 4.1100 1.1050 4.3000 1.1950 ;
      RECT 2.1250 0.4800 5.7150 0.5700 ;
      RECT 5.6250 0.5700 5.7150 1.5350 ;
      RECT 3.5500 1.0550 3.6400 1.4650 ;
      RECT 3.2750 0.9650 3.6400 1.0550 ;
      RECT 3.2750 0.5700 3.3650 0.9650 ;
      RECT 2.1250 0.5700 2.2150 1.3900 ;
      RECT 2.3700 0.4250 2.5400 0.4800 ;
      RECT 5.6100 1.6450 6.3200 1.7350 ;
      RECT 6.2300 1.4250 6.3200 1.6450 ;
      RECT 5.8150 0.6100 6.3200 0.7000 ;
      RECT 6.2300 0.4450 6.3200 0.6100 ;
      RECT 2.3800 1.8300 5.7000 1.9200 ;
      RECT 5.6100 1.7350 5.7000 1.8300 ;
      RECT 5.8150 0.7000 5.9050 1.6450 ;
      RECT 3.2350 1.4300 3.3250 1.8300 ;
      RECT 3.2350 1.2600 3.3700 1.4300 ;
  END
END M2DFFQ_X3M_A12TH

MACRO M2DFFQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.2450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.6900 ;
        RECT 2.7650 0.3200 2.9350 0.3800 ;
        RECT 3.3100 0.3200 3.4800 0.3800 ;
        RECT 6.6800 0.3200 6.8500 0.5050 ;
    END
  END VSS

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9800 1.5500 1.4050 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END D0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.2450 2.7200 ;
        RECT 0.3000 1.8800 0.5100 2.0800 ;
        RECT 1.6600 1.7350 1.7500 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3850 1.0500 5.9950 1.1500 ;
        RECT 5.3850 1.1500 5.4750 1.7300 ;
        RECT 5.9050 1.1500 5.9950 1.7150 ;
        RECT 5.3850 0.7000 5.4750 1.0500 ;
        RECT 5.9050 0.7000 5.9950 1.0500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8500 0.8350 6.9550 1.2600 ;
    END
    ANTENNAGATEAREA 0.0594 ;
  END CK

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4500 ;
    END
    ANTENNAGATEAREA 0.1044 ;
  END S0

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8000 0.5500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 0.6400 0.6900 0.7300 1.5800 ;
      RECT 0.6000 0.5200 0.7300 0.6900 ;
      RECT 0.0550 1.7000 0.9100 1.7900 ;
      RECT 0.8200 1.1050 0.9100 1.7000 ;
      RECT 0.2550 0.8900 0.3450 1.7000 ;
      RECT 0.0950 0.8000 0.3450 0.8900 ;
      RECT 0.0950 0.4800 0.1850 0.8000 ;
      RECT 1.2600 0.7600 1.3500 1.6750 ;
      RECT 1.0950 0.6700 1.3500 0.7600 ;
      RECT 1.6600 1.0600 1.8500 1.1500 ;
      RECT 1.7600 0.5700 1.8500 1.0600 ;
      RECT 0.8900 0.4800 1.8500 0.5700 ;
      RECT 0.8900 0.5700 0.9800 0.8650 ;
      RECT 0.8900 0.8650 1.0900 0.9550 ;
      RECT 1.0000 0.9550 1.0900 1.6750 ;
      RECT 1.9400 0.4800 2.0300 1.8900 ;
      RECT 2.2000 1.5900 2.2900 1.9250 ;
      RECT 2.2000 1.5000 2.3950 1.5900 ;
      RECT 2.3050 0.7550 2.3950 1.5000 ;
      RECT 2.3050 0.6650 2.9650 0.7550 ;
      RECT 2.8750 0.7550 2.9650 1.1750 ;
      RECT 2.6100 1.5700 3.6850 1.6600 ;
      RECT 3.5950 1.4750 3.6850 1.5700 ;
      RECT 2.6100 1.1150 2.7000 1.5700 ;
      RECT 3.0550 1.1050 3.1450 1.5700 ;
      RECT 3.0550 1.0150 3.1800 1.1050 ;
      RECT 3.0900 0.7550 3.1800 1.0150 ;
      RECT 3.0900 0.6650 3.7100 0.7550 ;
      RECT 3.6200 0.7550 3.7100 0.8750 ;
      RECT 4.4750 1.6250 5.0250 1.7150 ;
      RECT 4.4750 1.0400 4.5650 1.6250 ;
      RECT 4.9350 0.9500 5.0250 1.6250 ;
      RECT 4.8350 0.8600 5.0250 0.9500 ;
      RECT 3.9800 1.6500 4.3850 1.7400 ;
      RECT 4.2950 0.7500 4.3850 1.6500 ;
      RECT 4.0000 0.6600 5.2350 0.7500 ;
      RECT 4.0000 0.7500 4.0900 0.8450 ;
      RECT 4.6550 0.7500 4.7450 1.1050 ;
      RECT 5.1450 0.7500 5.2350 1.2250 ;
      RECT 4.6550 1.1050 4.8450 1.1950 ;
      RECT 2.1250 0.4800 6.5050 0.5700 ;
      RECT 6.4150 0.5700 6.5050 1.5750 ;
      RECT 4.0950 1.1500 4.1850 1.5600 ;
      RECT 3.4450 1.0600 4.1850 1.1500 ;
      RECT 3.4450 0.9150 3.5350 1.0600 ;
      RECT 3.8200 0.5700 3.9100 1.0600 ;
      RECT 2.1250 0.5700 2.2150 1.3900 ;
      RECT 2.3700 0.4500 2.5400 0.4800 ;
      RECT 6.4000 1.6900 7.1200 1.7800 ;
      RECT 7.0300 1.4450 7.1200 1.6900 ;
      RECT 6.6050 0.6100 7.1200 0.7000 ;
      RECT 7.0300 0.4750 7.1200 0.6100 ;
      RECT 6.6050 0.7000 6.6950 1.6900 ;
      RECT 2.3800 1.8300 6.4900 1.9200 ;
      RECT 6.4000 1.7800 6.4900 1.8300 ;
      RECT 3.7750 1.3400 3.8650 1.8300 ;
      RECT 3.4250 1.2500 3.8650 1.3400 ;
  END
END M2DFFQ_X4M_A12TH

MACRO M2SDFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.3350 0.3200 0.5050 0.6750 ;
        RECT 2.6250 0.3200 2.7950 0.4850 ;
        RECT 3.0650 0.3200 3.1750 0.4500 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8400 0.5950 1.3600 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8100 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0555 ;
  END S0

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5800 1.0500 3.0000 1.1500 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END SE

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8450 1.5500 1.2650 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D0

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2400 0.8350 7.3550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.8650 6.5500 1.4500 ;
        RECT 6.4500 1.4500 6.6400 1.5500 ;
        RECT 6.4500 0.7650 6.6750 0.8650 ;
        RECT 6.5400 1.5500 6.6400 1.6950 ;
    END
    ANTENNADIFFAREA 0.1304 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.4500 2.8700 1.5500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 2.5800 1.8450 2.7500 2.0800 ;
        RECT 0.3950 1.7000 0.4950 2.0800 ;
        RECT 3.1550 1.5050 3.2750 2.0800 ;
        RECT 1.5550 1.4950 1.6550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 5.4950 1.5250 6.3100 1.6150 ;
      RECT 5.4950 0.9650 5.5850 1.5250 ;
      RECT 6.2200 0.9500 6.3100 1.5250 ;
      RECT 5.9750 0.8600 6.3100 0.9500 ;
      RECT 3.6350 0.4800 6.8650 0.5700 ;
      RECT 6.7750 0.5700 6.8650 1.6550 ;
      RECT 4.9300 1.3000 5.1350 1.3900 ;
      RECT 4.9300 0.5700 5.0200 1.3000 ;
      RECT 3.6350 0.5700 3.7250 1.4350 ;
      RECT 3.8900 0.4350 4.0600 0.4800 ;
      RECT 6.9600 1.5000 7.5200 1.5900 ;
      RECT 7.4300 1.5900 7.5200 1.6700 ;
      RECT 6.9600 0.6100 7.5200 0.7000 ;
      RECT 7.4300 0.5300 7.5200 0.6100 ;
      RECT 3.8050 1.8200 7.0500 1.9100 ;
      RECT 6.9600 1.5900 7.0500 1.8200 ;
      RECT 6.9600 0.7000 7.0500 1.5000 ;
      RECT 0.7800 0.7300 0.8800 1.7150 ;
      RECT 0.6350 0.6400 0.8800 0.7300 ;
      RECT 0.8750 1.9150 1.0850 1.9650 ;
      RECT 0.5950 1.8250 1.0850 1.9150 ;
      RECT 0.5950 1.5900 0.6850 1.8250 ;
      RECT 0.0500 1.5000 0.6850 1.5900 ;
      RECT 0.0500 1.5900 0.1700 1.7300 ;
      RECT 0.0500 0.7300 0.1400 1.5000 ;
      RECT 0.0500 0.5600 0.2000 0.7300 ;
      RECT 1.3000 1.4850 1.3900 1.7000 ;
      RECT 1.1850 1.3950 1.3900 1.4850 ;
      RECT 1.1850 0.7500 1.2750 1.3950 ;
      RECT 1.1850 0.6600 1.3600 0.7500 ;
      RECT 0.9700 0.4800 1.9000 0.5700 ;
      RECT 1.8100 0.5700 1.9000 1.9450 ;
      RECT 0.9700 1.6050 1.1900 1.6950 ;
      RECT 0.9700 0.5700 1.0600 1.6050 ;
      RECT 2.8950 1.7500 2.9850 1.9600 ;
      RECT 2.2500 1.6600 2.9850 1.7500 ;
      RECT 2.2500 0.8600 3.0850 0.9500 ;
      RECT 2.9950 0.7600 3.0850 0.8600 ;
      RECT 2.2500 0.9500 2.3400 1.6600 ;
      RECT 2.0700 0.5750 3.3400 0.6650 ;
      RECT 3.2500 0.6650 3.3400 1.3600 ;
      RECT 2.0700 0.6650 2.1600 1.9250 ;
      RECT 3.4500 0.6050 3.5400 1.6950 ;
      RECT 3.6900 1.5550 3.9050 1.6450 ;
      RECT 3.8150 0.7700 3.9050 1.5550 ;
      RECT 3.8150 0.6800 4.5800 0.7700 ;
      RECT 4.4900 0.7700 4.5800 1.2950 ;
      RECT 4.1500 1.5250 4.7600 1.6150 ;
      RECT 4.1500 1.1100 4.2400 1.5250 ;
      RECT 4.6700 0.7700 4.7600 1.5250 ;
      RECT 4.6700 0.6800 4.8400 0.7700 ;
      RECT 4.8700 1.5550 5.3450 1.6450 ;
      RECT 5.2550 0.7700 5.3450 1.5550 ;
      RECT 5.1100 0.6800 5.8300 0.7700 ;
      RECT 5.7400 0.7700 5.8300 1.1100 ;
      RECT 5.7400 1.1100 5.9600 1.2000 ;
      RECT 5.8700 1.2000 5.9600 1.3200 ;
  END
END M2SDFFQN_X0P5M_A12TH

MACRO LATNRPQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6450 ;
        RECT 0.8450 0.3200 1.0150 0.5600 ;
        RECT 1.4300 0.3200 1.5200 0.6150 ;
        RECT 2.7300 0.3200 2.9000 0.4500 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.7100 2.0100 2.8000 2.0800 ;
        RECT 0.3400 1.7900 0.4300 2.0800 ;
        RECT 0.8600 1.7900 0.9500 2.0800 ;
        RECT 1.5500 1.5550 1.6400 2.0800 ;
    END
  END VDD

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.0800 1.1500 ;
        RECT 0.8100 0.8000 0.9100 1.0500 ;
    END
    ANTENNAGATEAREA 0.0774 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6450 1.0000 2.7500 1.4850 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.3700 2.3500 1.8200 ;
        RECT 2.2500 1.8200 2.7500 1.9200 ;
        RECT 2.0350 1.2700 2.3500 1.3700 ;
        RECT 2.6500 1.6650 2.7500 1.8200 ;
        RECT 2.0350 1.0600 2.1350 1.2700 ;
        RECT 2.6500 1.5750 2.9650 1.6650 ;
        RECT 1.9200 0.9700 2.1350 1.0600 ;
        RECT 2.8650 1.1700 2.9650 1.5750 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 0.6950 1.5500 ;
        RECT 0.0750 1.5500 0.1750 1.8600 ;
        RECT 0.5950 1.5500 0.6950 1.8600 ;
        RECT 0.0750 0.9500 0.1750 1.4500 ;
        RECT 0.0750 0.8500 0.6950 0.9500 ;
        RECT 0.5950 0.5300 0.6950 0.8500 ;
        RECT 0.0750 0.5150 0.1750 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN
  OBS
    LAYER M1 ;
      RECT 0.6100 1.2600 1.6500 1.3500 ;
      RECT 1.5600 1.3500 1.6500 1.4450 ;
      RECT 0.6100 1.1800 0.7000 1.2600 ;
      RECT 0.2850 1.0900 0.7000 1.1800 ;
      RECT 1.3200 1.3500 1.4100 1.7000 ;
      RECT 1.1700 0.4100 1.2600 1.2600 ;
      RECT 2.0700 1.5700 2.1600 1.9400 ;
      RECT 1.7400 1.4800 2.1600 1.5700 ;
      RECT 1.7400 0.4850 2.1600 0.5750 ;
      RECT 1.7400 1.1450 1.8300 1.4800 ;
      RECT 1.3500 1.0550 1.8300 1.1450 ;
      RECT 1.7400 0.5750 1.8300 1.0550 ;
      RECT 1.3500 0.9350 1.4400 1.0550 ;
      RECT 2.4400 0.7400 2.5300 1.7100 ;
      RECT 3.0300 1.7550 3.1450 1.9900 ;
      RECT 3.0550 0.6300 3.1450 1.7550 ;
      RECT 2.2500 0.5400 3.1450 0.6300 ;
      RECT 3.0300 0.4400 3.1450 0.5400 ;
      RECT 2.2500 0.6300 2.3400 1.1600 ;
  END
END LATNRPQN_X3M_A12TH

MACRO LATNRPQN_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.4150 0.3200 0.5850 0.3600 ;
        RECT 1.7650 0.3200 1.8550 0.6200 ;
        RECT 2.2850 0.3200 2.3750 0.6200 ;
        RECT 2.5900 0.3200 2.6800 0.6200 ;
        RECT 3.1100 0.3200 3.2000 0.6550 ;
        RECT 3.6300 0.3200 3.7200 0.6600 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.6200 1.1800 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.6500 1.0050 1.7500 ;
        RECT 0.4000 1.5700 0.5000 1.6500 ;
        RECT 0.9150 1.4350 1.0050 1.6500 ;
        RECT 0.2600 1.4800 0.5000 1.5700 ;
        RECT 0.9150 1.3450 1.2700 1.4350 ;
        RECT 0.2600 1.0900 0.3600 1.4800 ;
        RECT 1.1800 0.8750 1.2700 1.3450 ;
    END
    ANTENNAGATEAREA 0.1014 ;
  END GN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8200 1.0500 2.5600 1.1500 ;
        RECT 2.4700 1.1500 2.5600 1.2600 ;
        RECT 1.8200 0.9100 1.9150 1.0500 ;
    END
    ANTENNAGATEAREA 0.1272 ;
  END R

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.2500 3.5850 1.3500 ;
        RECT 2.8500 1.3500 2.9400 1.7200 ;
        RECT 3.3700 1.3500 3.4600 1.7200 ;
        RECT 3.4950 0.9800 3.5850 1.2500 ;
        RECT 2.8500 0.8900 3.5850 0.9800 ;
        RECT 2.8500 0.5500 2.9400 0.8900 ;
        RECT 3.3700 0.5500 3.4600 0.8900 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.4300 1.8950 0.6000 2.0800 ;
        RECT 1.6550 1.8400 1.7450 2.0800 ;
        RECT 2.5900 1.7700 2.6800 2.0800 ;
        RECT 3.1100 1.7700 3.2000 2.0800 ;
        RECT 3.6300 1.7700 3.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7300 0.6700 0.8200 1.5150 ;
      RECT 0.0800 0.4800 1.0200 0.5700 ;
      RECT 0.9300 0.5700 1.0200 1.2550 ;
      RECT 0.0800 0.5700 0.1700 1.7400 ;
      RECT 0.0800 0.4100 0.1700 0.4800 ;
      RECT 1.3600 1.2400 2.3400 1.3300 ;
      RECT 1.0950 1.6300 1.1850 1.9500 ;
      RECT 1.0950 1.5400 1.4500 1.6300 ;
      RECT 1.3600 1.3300 1.4500 1.5400 ;
      RECT 1.3600 0.7600 1.4500 1.2400 ;
      RECT 1.1100 0.6700 1.4500 0.7600 ;
      RECT 1.1100 0.5300 1.2000 0.6700 ;
      RECT 2.6500 1.0700 3.3850 1.1600 ;
      RECT 1.6200 0.8200 1.7100 1.0400 ;
      RECT 1.5400 1.0400 1.7100 1.1300 ;
      RECT 2.1150 1.5100 2.2050 1.8800 ;
      RECT 2.0250 0.4300 2.1150 0.7300 ;
      RECT 2.1150 1.4200 2.7400 1.5100 ;
      RECT 2.6500 1.1600 2.7400 1.4200 ;
      RECT 2.6500 0.8200 2.7400 1.0700 ;
      RECT 1.6200 0.7300 2.7400 0.8200 ;
  END
END LATNRPQN_X4M_A12TH

MACRO LATNRQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3600 0.3200 0.5300 0.4850 ;
        RECT 0.8550 0.3200 1.0250 0.4950 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.8100 2.3500 0.9400 ;
        RECT 2.1550 0.9400 2.3500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0350 0.9500 1.6400 ;
        RECT 0.8500 1.6400 2.4200 1.7400 ;
        RECT 2.3200 1.5500 2.4200 1.6400 ;
        RECT 2.3200 1.4500 2.6100 1.5500 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END RN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 1.3850 2.0100 1.5550 2.0800 ;
    END
  END VDD

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9400 2.7650 1.2500 ;
        RECT 1.8000 1.2500 2.7650 1.3500 ;
        RECT 1.8000 1.1800 1.9000 1.2500 ;
    END
    ANTENNAGATEAREA 0.0471 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5550 0.1700 1.7050 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q
  OBS
    LAYER M1 ;
      RECT 0.6500 0.8200 1.3300 0.9100 ;
      RECT 1.2400 0.9100 1.3300 1.2600 ;
      RECT 0.6500 0.9100 0.7400 1.4700 ;
      RECT 0.4700 1.8300 1.8500 1.9200 ;
      RECT 0.4700 0.5850 1.6850 0.6750 ;
      RECT 1.5950 0.4300 1.6850 0.5850 ;
      RECT 0.4700 1.1900 0.5600 1.8300 ;
      RECT 0.2650 1.0200 0.5600 1.1900 ;
      RECT 0.4700 0.6750 0.5600 1.0200 ;
      RECT 1.6200 1.4500 2.2000 1.5400 ;
      RECT 1.6200 0.9700 2.0650 1.0600 ;
      RECT 1.9750 0.6600 2.0650 0.9700 ;
      RECT 1.6200 1.0600 1.7100 1.4500 ;
      RECT 2.8100 1.6500 2.9450 1.8600 ;
      RECT 2.8550 0.7000 2.9450 1.6500 ;
      RECT 2.8050 0.5700 2.9450 0.7000 ;
      RECT 1.7750 0.4800 2.9450 0.5700 ;
      RECT 1.4200 0.8800 1.5100 1.4300 ;
      RECT 1.0500 1.4300 1.5100 1.5200 ;
      RECT 1.0500 1.3300 1.1400 1.4300 ;
      RECT 1.7750 0.5700 1.8650 0.7900 ;
      RECT 1.4200 0.7900 1.8650 0.8800 ;
  END
END LATNRQ_X0P5M_A12TH

MACRO LATNRQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.2850 0.3200 0.7150 0.3950 ;
        RECT 0.8500 0.3200 1.0200 0.4950 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.8100 2.3500 0.9400 ;
        RECT 2.1550 0.9400 2.3500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.8950 2.7650 1.2500 ;
        RECT 1.8000 1.2500 2.7650 1.3500 ;
        RECT 1.8000 1.1800 1.9100 1.2500 ;
    END
    ANTENNAGATEAREA 0.0792 ;
  END GN

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.0100 0.9500 1.6400 ;
        RECT 0.8500 1.6400 2.4200 1.7400 ;
        RECT 2.3200 1.5500 2.4200 1.6400 ;
        RECT 2.3200 1.4500 2.6100 1.5500 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END RN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5300 0.1700 1.7200 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 1.3700 2.0450 1.5400 2.0800 ;
        RECT 2.2750 1.8450 2.4450 2.0800 ;
        RECT 2.5650 1.7500 2.6650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6500 0.8000 1.3300 0.8900 ;
      RECT 1.2400 0.8900 1.3300 1.1600 ;
      RECT 0.6500 0.8900 0.7400 1.4900 ;
      RECT 0.4600 1.8300 1.8500 1.9200 ;
      RECT 0.8200 1.9200 1.0250 1.9800 ;
      RECT 0.4600 0.5850 1.6850 0.6750 ;
      RECT 1.5950 0.4300 1.6850 0.5850 ;
      RECT 0.4600 1.2100 0.5550 1.8300 ;
      RECT 0.2600 1.0400 0.5550 1.2100 ;
      RECT 0.4600 0.6750 0.5550 1.0400 ;
      RECT 1.6200 1.4500 2.2000 1.5400 ;
      RECT 1.6200 0.9700 2.0650 1.0600 ;
      RECT 1.9750 0.6600 2.0650 0.9700 ;
      RECT 1.6200 1.0600 1.7100 1.4500 ;
      RECT 2.8300 1.5800 2.9500 1.9700 ;
      RECT 2.8600 0.7300 2.9500 1.5800 ;
      RECT 2.8300 0.5700 2.9500 0.7300 ;
      RECT 1.7750 0.4800 2.9500 0.5700 ;
      RECT 1.4200 0.8800 1.5100 1.4300 ;
      RECT 1.0450 1.4300 1.5100 1.5200 ;
      RECT 1.0450 1.3400 1.1400 1.4300 ;
      RECT 1.7750 0.5700 1.8650 0.7900 ;
      RECT 1.4200 0.7900 1.8650 0.8800 ;
  END
END LATNRQ_X1M_A12TH

MACRO LATNRQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3750 0.3200 0.4650 0.6100 ;
        RECT 0.8450 0.3200 1.2450 0.3550 ;
        RECT 2.8350 0.3200 3.0450 0.3900 ;
    END
  END VSS

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.5800 1.3500 0.9750 ;
        RECT 0.9650 0.9750 1.3500 1.0750 ;
        RECT 1.2500 0.4800 3.1400 0.5800 ;
        RECT 3.0400 0.5800 3.1400 1.1400 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END RN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4100 1.2500 2.7500 1.3500 ;
        RECT 2.6500 1.1000 2.7500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 1.4500 3.1200 1.5500 ;
        RECT 2.2100 1.2800 2.3000 1.4500 ;
        RECT 2.0150 1.1900 2.3000 1.2800 ;
    END
    ANTENNAGATEAREA 0.0942 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 0.8500 0.7300 0.9500 ;
        RECT 0.2600 0.9500 0.3600 1.3350 ;
        RECT 0.6300 0.4850 0.7300 0.8500 ;
        RECT 0.2600 1.3350 0.6950 1.4350 ;
        RECT 0.5950 1.4350 0.6950 1.5500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 2.5100 1.8800 2.6800 2.0800 ;
        RECT 2.9300 1.8750 3.1000 2.0800 ;
        RECT 0.8600 1.8400 0.9500 2.0800 ;
        RECT 0.3400 1.8200 0.4300 2.0800 ;
        RECT 1.1200 1.8200 1.2100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0700 1.6400 1.3650 1.7300 ;
      RECT 1.2750 1.4500 1.3650 1.6400 ;
      RECT 1.2750 1.3600 1.4850 1.4500 ;
      RECT 0.0700 0.7350 0.1700 1.6400 ;
      RECT 1.8300 1.6400 1.9200 1.7400 ;
      RECT 1.6350 1.5500 1.9200 1.6400 ;
      RECT 1.6350 1.2550 1.7250 1.5500 ;
      RECT 0.7400 1.1650 1.7250 1.2550 ;
      RECT 1.6350 0.9200 1.7250 1.1650 ;
      RECT 1.6350 0.8300 1.9550 0.9200 ;
      RECT 1.6350 0.7350 1.7250 0.8300 ;
      RECT 1.8650 0.6900 1.9550 0.8300 ;
      RECT 0.7400 1.1500 0.8300 1.1650 ;
      RECT 0.4500 1.0600 0.8300 1.1500 ;
      RECT 1.0950 1.2550 1.1850 1.5000 ;
      RECT 2.0300 1.6500 2.2200 1.7400 ;
      RECT 2.0450 0.7100 2.3450 0.8000 ;
      RECT 1.8150 1.1000 1.9050 1.3700 ;
      RECT 2.0300 1.4600 2.1200 1.6500 ;
      RECT 1.8150 1.3700 2.1200 1.4600 ;
      RECT 1.8150 1.0100 2.1350 1.1000 ;
      RECT 2.0450 0.8000 2.1350 1.0100 ;
      RECT 2.3300 1.6800 3.3200 1.7700 ;
      RECT 3.2300 1.7700 3.3200 1.9700 ;
      RECT 3.2300 1.3400 3.3200 1.6800 ;
      RECT 2.8600 1.2500 3.3200 1.3400 ;
      RECT 3.2300 0.4600 3.3200 1.2500 ;
      RECT 2.8600 0.9000 2.9500 1.2500 ;
      RECT 2.4550 0.8100 2.9500 0.9000 ;
      RECT 1.4550 1.8300 2.4200 1.9200 ;
      RECT 2.3300 1.7700 2.4200 1.8300 ;
      RECT 1.4550 1.5600 1.5450 1.8300 ;
      RECT 2.4550 0.9000 2.5450 0.9400 ;
      RECT 2.2450 0.9400 2.5450 1.0500 ;
  END
END LATNRQ_X2M_A12TH

MACRO LATNRQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6850 ;
        RECT 0.8600 0.3200 0.9500 0.4650 ;
        RECT 1.2050 0.3200 1.3750 0.4800 ;
        RECT 3.1050 0.3200 3.1950 0.4250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.8600 1.9900 0.9500 2.0800 ;
        RECT 1.8900 1.9900 2.0600 2.0800 ;
        RECT 2.8700 1.9750 2.9600 2.0800 ;
        RECT 0.3400 1.7700 0.4300 2.0800 ;
        RECT 3.1350 1.6450 3.2250 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6100 0.8500 2.8700 0.9550 ;
        RECT 2.6800 0.9550 2.8700 1.0750 ;
    END
    ANTENNAGATEAREA 0.0966 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0100 1.0450 3.3000 1.1500 ;
        RECT 3.0100 1.1500 3.1000 1.1650 ;
        RECT 3.2100 1.1500 3.3000 1.2350 ;
        RECT 2.4800 1.1650 3.1000 1.2550 ;
        RECT 2.4800 1.2550 2.5700 1.3300 ;
        RECT 2.4800 1.1600 2.5700 1.1650 ;
    END
    ANTENNAGATEAREA 0.1005 ;
  END GN

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.4750 2.9500 1.7500 ;
        RECT 2.3700 1.7500 2.9500 1.8400 ;
        RECT 2.8500 1.3750 3.1600 1.4750 ;
        RECT 2.3700 1.7200 2.4600 1.7500 ;
        RECT 1.3400 1.6200 2.4600 1.7200 ;
        RECT 1.3400 1.1950 1.4300 1.6200 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END RN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 0.6950 1.5500 ;
        RECT 0.0750 1.5500 0.1750 1.8800 ;
        RECT 0.5950 1.5500 0.6950 1.8800 ;
        RECT 0.0750 0.9800 0.1700 1.4500 ;
        RECT 0.0750 0.8800 0.6950 0.9800 ;
        RECT 0.0750 0.5400 0.1750 0.8800 ;
        RECT 0.5950 0.5400 0.6950 0.8800 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q
  OBS
    LAYER M1 ;
      RECT 1.1450 0.9950 1.5800 1.0850 ;
      RECT 1.4900 0.8750 1.5800 0.9950 ;
      RECT 1.1450 1.0850 1.2350 1.6700 ;
      RECT 1.1450 0.7900 1.2350 0.9950 ;
      RECT 2.1000 1.3150 2.1900 1.4300 ;
      RECT 1.8700 1.2250 2.1900 1.3150 ;
      RECT 1.8700 0.9600 1.9600 1.2250 ;
      RECT 1.2950 1.9000 1.3850 1.9900 ;
      RECT 0.8700 1.8100 2.2800 1.9000 ;
      RECT 2.1900 1.9000 2.2800 1.9900 ;
      RECT 0.8700 0.6000 2.0650 0.6900 ;
      RECT 1.9750 0.4100 2.0650 0.6000 ;
      RECT 0.8700 1.1800 0.9600 1.8100 ;
      RECT 0.3400 1.0900 0.9600 1.1800 ;
      RECT 0.8700 0.6900 0.9600 1.0900 ;
      RECT 2.5700 1.5300 2.6600 1.6550 ;
      RECT 2.3000 1.4400 2.6600 1.5300 ;
      RECT 2.4100 0.6600 2.6200 0.7600 ;
      RECT 2.3000 0.9600 2.5000 1.0500 ;
      RECT 2.4100 0.7600 2.5000 0.9600 ;
      RECT 2.3000 1.0500 2.3900 1.4400 ;
      RECT 2.2300 0.5500 3.4850 0.5700 ;
      RECT 2.9250 0.5700 3.4850 0.6400 ;
      RECT 3.3950 0.6400 3.4850 1.9450 ;
      RECT 1.5450 1.4400 1.7600 1.5300 ;
      RECT 1.6700 0.8700 1.7600 1.4400 ;
      RECT 1.6700 0.7800 2.3200 0.8700 ;
      RECT 2.1000 0.8700 2.1900 1.1350 ;
      RECT 2.2300 0.5700 2.3200 0.7800 ;
      RECT 2.2300 0.4800 3.0150 0.5500 ;
  END
END LATNRQ_X3M_A12TH

MACRO LATNSPQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3700 0.3200 0.5600 0.4600 ;
        RECT 1.8100 0.3200 2.0150 0.5300 ;
        RECT 2.4950 0.3200 2.7000 0.7600 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7800 0.7500 1.2100 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0650 0.5500 1.5000 ;
        RECT 0.4500 1.5000 0.9250 1.5900 ;
        RECT 0.8350 1.5900 0.9250 1.6100 ;
        RECT 0.8350 1.6100 1.8400 1.7100 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END S

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8100 1.2900 2.9500 1.5000 ;
        RECT 2.8500 0.9700 2.9500 1.2900 ;
        RECT 2.8100 0.7600 2.9500 0.9700 ;
    END
    ANTENNADIFFAREA 0.14175 ;
  END Q

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.5700 1.1500 1.2400 ;
        RECT 0.6500 0.4800 1.6200 0.5700 ;
        RECT 0.0900 0.5700 0.7400 0.6700 ;
        RECT 1.5300 0.5700 1.6200 0.8000 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END GN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.2900 1.8700 0.5050 2.0800 ;
        RECT 2.5550 1.5350 2.6450 2.0800 ;
        RECT 1.9400 1.5150 2.0300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8150 1.3200 0.9850 1.4100 ;
      RECT 0.8500 0.6600 0.9400 1.3200 ;
      RECT 0.6350 1.8100 1.4000 1.9000 ;
      RECT 0.6350 1.7800 0.7250 1.8100 ;
      RECT 0.0800 1.6800 0.7250 1.7800 ;
      RECT 0.0800 0.8000 0.1700 1.6800 ;
      RECT 1.2600 0.8900 2.0350 0.9800 ;
      RECT 1.9450 0.9800 2.0350 1.0800 ;
      RECT 1.9450 0.7350 2.0350 0.8900 ;
      RECT 1.9450 1.0800 2.4150 1.1700 ;
      RECT 1.9450 0.6450 2.2200 0.7350 ;
      RECT 2.1300 0.4100 2.2200 0.6450 ;
      RECT 1.0950 1.3500 1.3500 1.4400 ;
      RECT 1.2600 0.9800 1.3500 1.3500 ;
      RECT 1.2600 0.6600 1.3500 0.8900 ;
      RECT 1.4800 1.3150 2.6150 1.4050 ;
      RECT 1.4800 1.0700 1.5700 1.3150 ;
      RECT 2.5250 0.9400 2.6150 1.3150 ;
      RECT 2.1500 0.8500 2.6150 0.9400 ;
  END
END LATNSPQ_X0P5M_A12TH

MACRO LATNSPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3400 0.3200 0.5300 0.4600 ;
        RECT 1.7950 0.3200 2.0050 0.5200 ;
        RECT 2.5500 0.3200 2.6400 0.6850 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9900 2.9500 1.2900 ;
        RECT 2.8050 1.2900 2.9500 1.3900 ;
        RECT 2.8050 0.8900 2.9500 0.9900 ;
        RECT 2.8050 1.3900 2.9000 1.6850 ;
        RECT 2.8050 0.5800 2.9000 0.8900 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7800 0.7500 1.2000 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END D

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0650 0.5500 1.5000 ;
        RECT 0.4500 1.5000 0.9250 1.6000 ;
        RECT 0.8350 1.6000 0.9250 1.6100 ;
        RECT 0.8350 1.6100 1.8400 1.7100 ;
    END
    ANTENNAGATEAREA 0.0786 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 2.5500 1.7700 2.6400 2.0800 ;
        RECT 1.9400 1.5000 2.0300 2.0800 ;
    END
  END VDD

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.5700 1.1500 1.2300 ;
        RECT 0.0900 0.5500 1.6100 0.5700 ;
        RECT 0.0900 0.5700 0.7300 0.6500 ;
        RECT 1.5200 0.5700 1.6100 0.8000 ;
        RECT 0.6400 0.4800 1.6100 0.5500 ;
    END
    ANTENNAGATEAREA 0.0624 ;
  END GN
  OBS
    LAYER M1 ;
      RECT 0.7950 1.3200 0.9850 1.4100 ;
      RECT 0.8400 0.6600 0.9300 1.3200 ;
      RECT 0.0950 1.8100 1.4000 1.9000 ;
      RECT 0.0950 0.7800 0.1850 1.8100 ;
      RECT 1.2600 0.8900 2.0550 0.9800 ;
      RECT 1.9650 0.9800 2.0550 1.0800 ;
      RECT 1.9650 0.7350 2.0550 0.8900 ;
      RECT 1.9650 1.0800 2.4350 1.1700 ;
      RECT 1.9650 0.6450 2.2200 0.7350 ;
      RECT 2.1300 0.4100 2.2200 0.6450 ;
      RECT 1.0950 1.3700 1.3500 1.4600 ;
      RECT 1.2600 0.9800 1.3500 1.3700 ;
      RECT 1.2600 0.6600 1.3500 0.8900 ;
      RECT 1.4800 1.3200 2.6150 1.4100 ;
      RECT 1.4800 1.0700 1.5700 1.3200 ;
      RECT 2.5250 0.9400 2.6150 1.3200 ;
      RECT 2.1650 0.8500 2.6150 0.9400 ;
  END
END LATNSPQ_X1M_A12TH

MACRO LATNSPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3500 0.3200 0.5400 0.4600 ;
        RECT 1.7800 0.3200 1.9900 0.5300 ;
        RECT 2.5100 0.3200 2.6000 0.6900 ;
        RECT 3.0300 0.3200 3.1200 0.6850 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7700 0.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.5700 1.1500 1.2550 ;
        RECT 0.0950 0.5500 1.5950 0.5700 ;
        RECT 0.0950 0.5700 0.7400 0.6500 ;
        RECT 1.5050 0.5700 1.5950 0.8000 ;
        RECT 0.6500 0.4800 1.5950 0.5500 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9700 2.9500 1.2900 ;
        RECT 2.7700 1.2900 2.9500 1.3900 ;
        RECT 2.7700 0.8500 2.9500 0.9700 ;
        RECT 2.7700 1.3900 2.8600 1.7200 ;
        RECT 2.7700 0.5400 2.8600 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0650 0.5500 1.6000 ;
        RECT 0.4500 1.6000 1.8500 1.7000 ;
    END
    ANTENNAGATEAREA 0.0786 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.5100 1.7700 2.6000 2.0800 ;
        RECT 3.0300 1.7700 3.1200 2.0800 ;
        RECT 1.9400 1.5200 2.0300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8500 0.6600 0.9400 1.5000 ;
      RECT 0.0950 1.8100 1.4200 1.9000 ;
      RECT 0.0950 0.7600 0.1850 1.8100 ;
      RECT 1.2600 0.8900 2.0100 0.9800 ;
      RECT 1.9200 0.9800 2.0100 1.0800 ;
      RECT 1.9200 0.7350 2.0100 0.8900 ;
      RECT 1.9200 1.0800 2.4150 1.1700 ;
      RECT 1.9200 0.6450 2.2050 0.7350 ;
      RECT 2.1150 0.4100 2.2050 0.6450 ;
      RECT 1.0750 1.3700 1.3500 1.4600 ;
      RECT 1.2600 0.9800 1.3500 1.3700 ;
      RECT 1.2600 0.6600 1.3500 0.8900 ;
      RECT 1.5200 1.3200 2.6300 1.4100 ;
      RECT 1.5200 1.0700 1.6100 1.3200 ;
      RECT 2.5400 0.9400 2.6300 1.3200 ;
      RECT 2.1200 0.8500 2.6300 0.9400 ;
  END
END LATNSPQ_X2M_A12TH

MACRO LATNSPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3800 0.3200 0.5900 0.5000 ;
        RECT 1.0600 0.3200 1.1500 0.5000 ;
        RECT 2.2100 0.3200 2.3100 0.8000 ;
        RECT 3.2350 0.3200 3.3250 0.6850 ;
        RECT 3.7700 0.3200 3.8600 0.6850 ;
    END
  END VSS

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0250 0.5500 1.5000 ;
        RECT 0.4400 1.5000 2.5400 1.5900 ;
        RECT 2.4500 1.5900 2.5400 1.9300 ;
        RECT 1.2500 1.0250 1.3400 1.5000 ;
    END
    ANTENNAGATEAREA 0.1332 ;
  END S

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0100 0.9000 1.1900 ;
    END
    ANTENNAGATEAREA 0.1527 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.5700 1.9500 0.7900 ;
        RECT 1.4400 0.4800 1.9500 0.5700 ;
        RECT 1.4400 0.5700 1.5300 0.5900 ;
        RECT 0.1500 0.5900 1.5300 0.6900 ;
        RECT 0.1500 0.4100 0.2400 0.5900 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5050 1.0500 4.1250 1.1500 ;
        RECT 3.5050 1.1500 3.6050 1.7200 ;
        RECT 4.0250 1.1500 4.1250 1.7200 ;
        RECT 3.5050 0.5400 3.6050 1.0500 ;
        RECT 4.0250 0.5400 4.1250 1.0500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 3.2500 1.7700 3.3400 2.0800 ;
        RECT 3.7700 1.7700 3.8600 2.0800 ;
        RECT 2.6400 1.5000 2.8100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.7700 2.2400 1.8600 ;
      RECT 0.0800 0.7900 0.1700 1.7700 ;
      RECT 1.6400 0.8900 2.7150 0.9800 ;
      RECT 2.6250 0.9800 2.7150 1.0800 ;
      RECT 2.6250 0.6450 2.7150 0.8900 ;
      RECT 2.6250 1.0800 3.1550 1.1700 ;
      RECT 1.8800 1.3200 2.0850 1.4100 ;
      RECT 1.9950 0.9800 2.0850 1.3200 ;
      RECT 1.6400 0.6650 1.7300 0.8900 ;
      RECT 2.2900 1.3200 3.3550 1.4100 ;
      RECT 2.2900 1.0700 2.3800 1.3200 ;
      RECT 3.2650 0.9400 3.3550 1.3200 ;
      RECT 2.8250 0.8500 3.3550 0.9400 ;
      RECT 0.7150 0.8000 1.5400 0.8900 ;
      RECT 1.4500 0.8900 1.5400 1.3200 ;
      RECT 1.4500 1.3200 1.7700 1.4100 ;
      RECT 0.7400 1.3200 1.1400 1.4100 ;
      RECT 1.0500 0.8900 1.1400 1.3200 ;
  END
END LATNSPQ_X3M_A12TH

MACRO LATNSQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 1.1950 0.3200 1.2950 0.6050 ;
        RECT 0.3350 0.3200 0.4350 0.6900 ;
        RECT 2.2300 0.3200 2.4000 0.7800 ;
        RECT 0.9850 0.6050 1.2950 0.7050 ;
        RECT 0.9850 0.7050 1.0850 0.8850 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8400 0.5600 1.2600 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0700 1.0500 2.4900 1.1500 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.4650 1.7500 1.8200 ;
        RECT 1.6500 1.8200 2.2500 1.9200 ;
        RECT 1.4050 1.3650 1.7500 1.4650 ;
        RECT 2.1500 1.5500 2.2500 1.8200 ;
        RECT 1.4050 0.9800 1.5050 1.3650 ;
        RECT 2.1500 1.4500 2.5500 1.5500 ;
        RECT 2.4400 1.3350 2.5500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.4100 0.1700 1.8900 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.3500 1.7200 0.4500 2.0800 ;
        RECT 2.3400 1.6900 2.4400 2.0800 ;
        RECT 0.9500 1.6800 1.0500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6750 0.9950 1.1000 1.1650 ;
      RECT 0.7850 0.4250 1.0650 0.5150 ;
      RECT 0.6750 1.5900 0.7650 1.8900 ;
      RECT 0.2600 1.5000 0.7650 1.5900 ;
      RECT 0.6750 1.1650 0.7650 1.5000 ;
      RECT 0.7850 0.5150 0.8750 0.9950 ;
      RECT 0.2600 1.1100 0.3500 1.5000 ;
      RECT 1.4500 1.6450 1.5400 1.8600 ;
      RECT 1.2050 1.5550 1.5400 1.6450 ;
      RECT 1.2050 0.8000 1.6000 0.8900 ;
      RECT 1.5100 0.6650 1.6000 0.8000 ;
      RECT 1.2050 1.4300 1.2950 1.5550 ;
      RECT 0.8550 1.3300 1.2950 1.4300 ;
      RECT 1.2050 0.8900 1.2950 1.3300 ;
      RECT 1.8700 1.6400 2.0400 1.7300 ;
      RECT 1.8700 0.6900 1.9600 1.6400 ;
      RECT 2.5450 1.7400 2.7350 1.8500 ;
      RECT 2.6450 0.9600 2.7350 1.7400 ;
      RECT 2.0500 0.8700 2.7350 0.9600 ;
      RECT 2.6100 0.6450 2.7350 0.8700 ;
      RECT 2.0500 0.5800 2.1400 0.8700 ;
      RECT 1.6900 0.4900 2.1400 0.5800 ;
      RECT 1.6900 0.5800 1.7800 1.2550 ;
  END
END LATNSQN_X0P5M_A12TH

MACRO LATNSQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6950 ;
        RECT 1.1000 0.3200 1.2000 0.6900 ;
        RECT 2.3700 0.3200 2.4700 0.7000 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4700 0.8700 0.7500 0.9900 ;
        RECT 0.6500 0.6150 0.7500 0.8700 ;
    END
    ANTENNAGATEAREA 0.0558 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2450 1.0100 2.3500 1.2900 ;
        RECT 2.1400 1.2900 2.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.0400 2.5650 1.5700 ;
        RECT 2.1600 1.5700 2.5650 1.6700 ;
        RECT 2.1600 1.6700 2.2600 1.8200 ;
        RECT 1.7500 1.8200 2.2600 1.9200 ;
        RECT 1.7500 1.3700 1.8500 1.8200 ;
        RECT 1.4950 1.2700 1.8500 1.3700 ;
        RECT 1.4950 0.8700 1.5950 1.2700 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5150 0.1700 1.7000 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.3400 1.8000 0.4400 2.0800 ;
        RECT 0.9300 1.7900 1.0300 2.0800 ;
        RECT 2.3700 1.7800 2.4700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8650 0.9600 1.1900 1.0700 ;
      RECT 0.2600 1.0900 0.9550 1.1800 ;
      RECT 0.8650 1.0700 0.9550 1.0900 ;
      RECT 0.8650 0.4100 0.9550 0.9600 ;
      RECT 0.5500 1.8300 0.8050 1.9200 ;
      RECT 0.5500 1.1800 0.6400 1.8300 ;
      RECT 1.2950 1.8200 1.6550 1.9100 ;
      RECT 1.2950 0.6900 1.6500 0.7800 ;
      RECT 1.5600 0.4950 1.6500 0.6900 ;
      RECT 1.2950 1.3800 1.3850 1.8200 ;
      RECT 0.7600 1.2900 1.3850 1.3800 ;
      RECT 1.2950 0.7800 1.3850 1.2900 ;
      RECT 0.7600 1.3800 0.8500 1.6800 ;
      RECT 1.9600 0.6600 2.0500 1.7300 ;
      RECT 2.6300 1.7350 2.7450 1.9450 ;
      RECT 2.6550 0.9000 2.7450 1.7350 ;
      RECT 2.1900 0.8100 2.7450 0.9000 ;
      RECT 2.6300 0.5450 2.7450 0.8100 ;
      RECT 1.7550 0.5700 1.8500 1.1800 ;
      RECT 2.1900 0.5700 2.2800 0.8100 ;
      RECT 1.7550 0.4800 2.2800 0.5700 ;
  END
END LATNSQN_X1M_A12TH

MACRO LATNSQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.5000 0.3200 0.6700 0.5850 ;
        RECT 1.0300 0.3200 1.2000 0.5850 ;
        RECT 2.3300 0.3200 2.4300 0.6200 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.1150 2.3500 1.4200 ;
        RECT 2.1500 1.0050 2.3500 1.1150 ;
    END
    ANTENNAGATEAREA 0.0558 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.9900 0.5500 1.4100 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END SN

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.1950 2.5500 1.6500 ;
        RECT 2.1700 1.6500 2.5500 1.7500 ;
        RECT 2.1700 1.7500 2.2700 1.8200 ;
        RECT 1.7800 1.8200 2.2700 1.9200 ;
        RECT 1.7800 1.3500 1.8800 1.8200 ;
        RECT 1.5000 1.2500 1.8800 1.3500 ;
        RECT 1.5000 0.8550 1.6000 1.2500 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9600 1.1500 1.2850 ;
        RECT 0.8500 1.2850 1.1500 1.3850 ;
        RECT 0.7500 0.8600 1.1500 0.9600 ;
        RECT 0.8500 1.3850 0.9500 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.3650 1.8650 2.4650 2.0800 ;
        RECT 0.0750 1.8200 0.1750 2.0800 ;
        RECT 0.5950 1.8200 0.6950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6600 1.0900 0.9400 1.1900 ;
      RECT 0.0800 1.6400 0.7500 1.7300 ;
      RECT 0.6600 1.1900 0.7500 1.6400 ;
      RECT 0.3400 1.7300 0.4300 1.9900 ;
      RECT 0.0800 0.5400 0.1700 1.6400 ;
      RECT 1.6000 1.5300 1.6900 1.6950 ;
      RECT 1.3000 1.4400 1.6900 1.5300 ;
      RECT 0.2650 0.6750 1.7000 0.7650 ;
      RECT 1.6100 0.4300 1.7000 0.6750 ;
      RECT 1.3000 0.7650 1.3900 1.4400 ;
      RECT 0.2650 0.7650 0.3550 1.5300 ;
      RECT 1.9700 0.6800 2.0600 1.7100 ;
      RECT 2.6100 1.8200 2.7300 1.9900 ;
      RECT 2.6400 0.8200 2.7300 1.8200 ;
      RECT 2.1500 0.7300 2.7300 0.8200 ;
      RECT 2.6300 0.5450 2.7300 0.7300 ;
      RECT 1.7900 0.5700 1.8800 1.1400 ;
      RECT 2.1500 0.5700 2.2400 0.7300 ;
      RECT 1.7900 0.4800 2.2400 0.5700 ;
  END
END LATNSQN_X2M_A12TH

MACRO LATNSQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.5000 0.3200 0.6700 0.5850 ;
        RECT 1.0300 0.3200 1.2000 0.5850 ;
        RECT 1.5700 0.3200 1.7400 0.5850 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.9900 0.5500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6350 0.9550 2.7500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9750 2.9550 1.6200 ;
        RECT 2.6500 1.6200 2.9550 1.7200 ;
        RECT 2.6500 1.7200 2.7500 1.8200 ;
        RECT 2.2650 1.8200 2.7500 1.9200 ;
        RECT 2.2650 1.3500 2.3650 1.8200 ;
        RECT 2.0150 1.2500 2.3650 1.3500 ;
        RECT 2.0150 0.8550 2.1150 1.2500 ;
    END
    ANTENNAGATEAREA 0.0816 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9600 1.5500 1.2850 ;
        RECT 0.8550 1.2850 1.5500 1.3850 ;
        RECT 0.7500 0.8600 1.5500 0.9600 ;
        RECT 0.8550 1.3850 0.9550 1.7200 ;
        RECT 1.3750 1.3850 1.4750 1.7150 ;
    END
    ANTENNADIFFAREA 0.602875 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.6850 2.0150 2.8950 2.0800 ;
        RECT 0.0750 1.8200 0.1750 2.0800 ;
        RECT 0.5950 1.8200 0.6950 2.0800 ;
        RECT 1.1150 1.7700 1.2150 2.0800 ;
        RECT 1.6250 1.4800 1.7250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6600 1.0900 1.2750 1.1900 ;
      RECT 0.3400 1.7300 0.4300 1.9900 ;
      RECT 0.0800 0.5400 0.1700 1.6400 ;
      RECT 0.0800 1.6400 0.7500 1.7300 ;
      RECT 0.6600 1.1900 0.7500 1.6400 ;
      RECT 2.0850 1.5300 2.1750 1.6950 ;
      RECT 1.8150 1.4400 2.1750 1.5300 ;
      RECT 0.2650 0.6750 2.1750 0.7650 ;
      RECT 2.0850 0.4450 2.1750 0.6750 ;
      RECT 1.8150 0.7650 1.9050 1.4400 ;
      RECT 0.2650 0.7650 0.3550 1.5300 ;
      RECT 2.4550 0.6800 2.5450 1.7100 ;
      RECT 3.0100 1.8150 3.1500 1.9900 ;
      RECT 3.0600 0.7750 3.1500 1.8150 ;
      RECT 3.0200 0.5700 3.1500 0.7750 ;
      RECT 2.2750 0.4800 3.1500 0.5700 ;
      RECT 2.2750 0.5700 2.3650 1.1350 ;
  END
END LATNSQN_X3M_A12TH

MACRO LATNSQN_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3250 0.3200 0.4950 0.4000 ;
        RECT 1.6550 0.3200 1.7550 0.6300 ;
        RECT 2.6450 0.3200 2.7450 0.6650 ;
        RECT 3.1650 0.3200 3.2650 0.6650 ;
    END
  END VSS

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.4550 0.9500 1.7900 ;
        RECT 0.4500 1.7900 0.9500 1.8800 ;
        RECT 0.8500 1.3550 1.1500 1.4550 ;
        RECT 0.4500 1.5150 0.5500 1.7900 ;
        RECT 1.0500 1.0350 1.1500 1.3550 ;
        RECT 0.2300 1.4150 0.5500 1.5150 ;
        RECT 1.0500 0.9350 1.3050 1.0350 ;
        RECT 0.2300 1.0000 0.3300 1.4150 ;
    END
    ANTENNAGATEAREA 0.1038 ;
  END GN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7700 0.5550 1.1850 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6750 1.0500 2.6350 1.1100 ;
        RECT 1.9450 1.1100 2.6350 1.1500 ;
        RECT 1.6750 1.0100 2.0350 1.0500 ;
        RECT 2.5350 1.1500 2.6350 1.2400 ;
    END
    ANTENNAGATEAREA 0.162 ;
  END SN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9100 1.2500 3.5250 1.3500 ;
        RECT 2.9100 1.3500 3.0100 1.7200 ;
        RECT 3.4250 1.3500 3.5250 1.7200 ;
        RECT 3.4250 0.9500 3.5250 1.2500 ;
        RECT 2.9100 0.8500 3.5250 0.9500 ;
        RECT 2.9100 0.5200 3.0100 0.8500 ;
        RECT 3.4250 0.5200 3.5250 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.3950 1.9900 0.4950 2.0800 ;
        RECT 1.6050 1.7700 1.7050 2.0800 ;
        RECT 2.1250 1.7700 2.2250 2.0800 ;
        RECT 2.6450 1.7700 2.7450 2.0800 ;
        RECT 3.1650 1.7700 3.2650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 0.4900 0.9300 0.5800 ;
      RECT 0.8400 0.5800 0.9300 1.2300 ;
      RECT 0.0500 1.6200 0.1700 1.9900 ;
      RECT 0.0500 0.5800 0.1400 1.6200 ;
      RECT 0.0500 0.4100 0.1700 0.4900 ;
      RECT 1.2450 1.2800 2.3800 1.2900 ;
      RECT 1.7550 1.2900 2.3800 1.3700 ;
      RECT 1.0400 1.6500 1.1300 1.9700 ;
      RECT 1.0400 1.5600 1.3350 1.6500 ;
      RECT 1.2450 1.2900 1.3350 1.5600 ;
      RECT 1.4600 0.7950 1.5500 1.2000 ;
      RECT 1.0400 0.7050 1.5500 0.7950 ;
      RECT 1.2450 1.2000 1.8450 1.2800 ;
      RECT 2.7300 1.0600 3.3150 1.1500 ;
      RECT 1.4450 1.3800 1.6550 1.4600 ;
      RECT 1.8700 1.5500 1.9600 1.9450 ;
      RECT 2.3900 1.5500 2.4800 1.9450 ;
      RECT 2.1300 0.5200 2.2200 0.8600 ;
      RECT 1.4450 1.4600 2.8200 1.5500 ;
      RECT 2.7300 1.1500 2.8200 1.4600 ;
      RECT 2.7300 0.9500 2.8200 1.0600 ;
      RECT 2.1300 0.8600 2.8200 0.9500 ;
      RECT 0.6600 0.6900 0.7500 1.6800 ;
  END
END LATNSQN_X4M_A12TH

MACRO LATQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 1.6800 0.3200 1.7700 0.7900 ;
        RECT 2.1700 0.3200 2.2600 0.9300 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.5800 0.5500 0.8450 ;
        RECT 0.4500 0.4800 1.1400 0.5800 ;
        RECT 0.2450 0.8450 0.5500 0.9500 ;
        RECT 1.0500 0.5800 1.1400 1.1650 ;
        RECT 1.0500 1.1650 1.3350 1.2550 ;
        RECT 1.2450 1.2550 1.3350 1.5350 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END G

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2100 0.6300 1.3900 ;
    END
    ANTENNAGATEAREA 0.0291 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4250 0.5250 2.5500 1.7200 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.3400 1.6650 0.4300 2.0800 ;
        RECT 1.6800 1.5950 1.7700 2.0800 ;
        RECT 2.1700 1.3150 2.2600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7400 1.6400 0.9300 1.7300 ;
      RECT 0.7400 0.7800 0.8300 1.6400 ;
      RECT 0.7400 0.6900 0.9500 0.7800 ;
      RECT 1.0400 1.9150 1.2100 1.9800 ;
      RECT 0.5400 1.8250 1.2100 1.9150 ;
      RECT 0.5400 1.5750 0.6300 1.8250 ;
      RECT 0.0500 1.4850 0.6300 1.5750 ;
      RECT 0.0500 1.5750 0.1750 1.8350 ;
      RECT 0.0500 0.7600 0.1400 1.4850 ;
      RECT 0.0500 0.5700 0.1750 0.7600 ;
      RECT 1.4250 1.0200 1.8500 1.1100 ;
      RECT 1.7600 0.9000 1.8500 1.0200 ;
      RECT 1.1400 1.6450 1.5150 1.7350 ;
      RECT 1.4250 1.1100 1.5150 1.6450 ;
      RECT 1.4250 0.8100 1.5150 1.0200 ;
      RECT 1.2300 0.7150 1.5150 0.8100 ;
      RECT 1.2300 0.6000 1.3200 0.7150 ;
      RECT 1.9400 1.0500 2.3050 1.1500 ;
      RECT 1.6050 1.3200 1.6950 1.4400 ;
      RECT 1.6050 1.2300 2.0300 1.3200 ;
      RECT 1.9400 1.3200 2.0300 1.8250 ;
      RECT 1.9400 1.1500 2.0300 1.2300 ;
      RECT 1.9400 0.6150 2.0300 1.0500 ;
  END
END LATQN_X0P5M_A12TH

MACRO LATQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 1.6300 0.3200 1.7200 0.7050 ;
        RECT 2.1700 0.3200 2.2600 0.6500 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9700 0.8500 1.2300 0.9500 ;
        RECT 1.1300 0.9500 1.2300 1.2600 ;
        RECT 0.9700 0.5800 1.0700 0.8500 ;
        RECT 1.1300 1.2600 1.3550 1.3600 ;
        RECT 0.4500 0.4800 1.0700 0.5800 ;
        RECT 0.4500 0.5800 0.5500 0.8550 ;
        RECT 0.2500 0.8550 0.5500 0.9500 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END G

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.1250 0.6100 1.3350 ;
        RECT 0.4500 1.3350 0.5500 1.5150 ;
    END
    ANTENNAGATEAREA 0.0372 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9350 2.5500 1.2950 ;
        RECT 2.4300 1.2950 2.5500 1.7250 ;
        RECT 2.4300 0.5050 2.5500 0.9350 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 2.1700 1.7700 2.2600 2.0800 ;
        RECT 1.6450 1.4200 1.7350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7200 0.7600 0.8100 1.6600 ;
      RECT 0.6600 0.6700 0.8600 0.7600 ;
      RECT 0.0550 1.7800 1.0100 1.8700 ;
      RECT 0.9200 1.1050 1.0100 1.7800 ;
      RECT 0.0550 1.5000 0.1700 1.7800 ;
      RECT 0.0550 0.7650 0.1450 1.5000 ;
      RECT 0.0550 0.5550 0.1700 0.7650 ;
      RECT 1.3300 1.0800 1.8400 1.1700 ;
      RECT 1.7500 1.1700 1.8400 1.2900 ;
      RECT 1.1000 1.5400 1.1900 1.6600 ;
      RECT 1.1000 1.4500 1.5550 1.5400 ;
      RECT 1.4650 1.1700 1.5550 1.4500 ;
      RECT 1.3300 0.7150 1.4200 1.0800 ;
      RECT 1.1650 0.6100 1.4200 0.7150 ;
      RECT 1.1650 0.5050 1.2550 0.6100 ;
      RECT 1.5300 0.8800 2.3400 0.9700 ;
      RECT 2.2500 0.9700 2.3400 1.2150 ;
      RECT 1.8650 1.4800 2.0400 1.7700 ;
      RECT 1.9500 0.9700 2.0400 1.4800 ;
      RECT 1.9050 0.4650 1.9950 0.8800 ;
      RECT 1.5300 0.7950 1.6300 0.8800 ;
  END
END LATQN_X1M_A12TH

MACRO LATQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3600 0.3200 0.5300 0.5100 ;
        RECT 0.8800 0.3200 1.0500 0.5100 ;
        RECT 2.2700 0.3200 2.3600 0.9000 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.2000 2.1600 1.5900 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.5700 1.7500 1.2000 ;
        RECT 1.6500 0.4800 2.1500 0.5700 ;
        RECT 2.0500 0.5700 2.1500 0.9900 ;
        RECT 2.0500 0.9900 2.5100 1.0900 ;
        RECT 2.4100 1.0900 2.5100 1.1600 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9050 0.9500 1.4900 ;
        RECT 0.6550 1.4900 0.9500 1.5900 ;
        RECT 0.6000 0.8050 0.9500 0.9050 ;
        RECT 0.6550 1.5900 0.7550 1.9200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.4000 1.7700 0.4900 2.0800 ;
        RECT 0.9200 1.7700 1.0100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.3000 0.6750 1.3900 ;
      RECT 0.5850 1.0150 0.6750 1.3000 ;
      RECT 0.0800 1.3900 0.1700 1.7200 ;
      RECT 0.0800 0.4900 0.1700 1.3000 ;
      RECT 1.4800 1.6000 1.5700 1.7000 ;
      RECT 1.1850 1.5100 1.5700 1.6000 ;
      RECT 1.1850 0.7150 1.2750 1.5100 ;
      RECT 1.1850 0.7050 1.5600 0.7150 ;
      RECT 0.2600 0.6150 1.5600 0.7050 ;
      RECT 1.4700 0.5250 1.5600 0.6150 ;
      RECT 0.2600 0.7050 0.3500 1.1900 ;
      RECT 1.8700 0.6800 1.9600 1.7200 ;
      RECT 1.6900 1.8300 2.7050 1.9200 ;
      RECT 2.6150 0.6800 2.7050 1.8300 ;
      RECT 1.3950 0.8600 1.4850 1.3300 ;
      RECT 1.6900 1.4200 1.7800 1.8300 ;
      RECT 1.3950 1.3300 1.7800 1.4200 ;
  END
END LATQN_X2M_A12TH

MACRO LATQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6850 ;
        RECT 1.7350 0.3200 1.8350 0.7650 ;
        RECT 2.2500 0.3200 2.3400 0.6850 ;
        RECT 2.7700 0.3200 2.8600 0.6850 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9500 0.3500 1.1950 ;
        RECT 0.2500 0.8500 0.6250 0.9500 ;
        RECT 0.5250 0.5800 0.6250 0.8500 ;
        RECT 0.5250 0.4800 1.0350 0.5800 ;
        RECT 0.9450 0.5800 1.0350 1.1850 ;
    END
    ANTENNAGATEAREA 0.0786 ;
  END G

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.3450 0.5500 1.5950 ;
        RECT 0.4500 1.2450 0.6400 1.3450 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5050 1.4500 3.1500 1.5500 ;
        RECT 2.5050 1.5500 2.6050 1.8800 ;
        RECT 3.0250 1.5500 3.1500 1.8800 ;
        RECT 3.0500 0.9500 3.1500 1.4500 ;
        RECT 2.5100 0.8500 3.1500 0.9500 ;
        RECT 2.5100 0.5200 2.6000 0.8500 ;
        RECT 3.0300 0.5200 3.1500 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3350 1.9400 0.4350 2.0800 ;
        RECT 1.7400 1.7700 1.8300 2.0800 ;
        RECT 2.2500 1.7700 2.3400 2.0800 ;
        RECT 2.7700 1.7700 2.8600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7350 0.6800 0.8250 1.6900 ;
      RECT 0.5200 1.8100 1.0300 1.9000 ;
      RECT 0.9400 1.3800 1.0300 1.8100 ;
      RECT 0.9400 1.2900 1.3350 1.3800 ;
      RECT 1.2450 0.8200 1.3350 1.2900 ;
      RECT 0.0650 1.7000 0.6100 1.7900 ;
      RECT 0.5200 1.7900 0.6100 1.8100 ;
      RECT 0.0650 1.7900 0.1700 1.9100 ;
      RECT 0.0650 0.7150 0.1550 1.7000 ;
      RECT 0.0650 0.5050 0.2100 0.7150 ;
      RECT 1.4450 0.9100 1.9450 1.0100 ;
      RECT 1.1400 1.5700 1.2300 1.8700 ;
      RECT 1.1400 1.4800 1.5350 1.5700 ;
      RECT 1.4450 1.0100 1.5350 1.4800 ;
      RECT 1.4450 0.7100 1.5350 0.9100 ;
      RECT 1.1250 0.6200 1.5350 0.7100 ;
      RECT 1.1250 0.5000 1.2350 0.6200 ;
      RECT 2.0700 1.0900 2.8300 1.1800 ;
      RECT 1.6250 1.1200 1.7150 1.2400 ;
      RECT 2.0000 1.3300 2.0900 1.7950 ;
      RECT 1.6250 1.2400 2.1600 1.3300 ;
      RECT 2.0700 1.1800 2.1600 1.2400 ;
      RECT 2.0700 0.8200 2.1600 1.0900 ;
      RECT 2.0000 0.7300 2.1600 0.8200 ;
      RECT 2.0000 0.4400 2.0900 0.7300 ;
  END
END LATQN_X3M_A12TH

MACRO LATQN_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 1.6800 0.3200 1.7700 0.6300 ;
        RECT 2.1850 0.3200 2.2850 0.6650 ;
        RECT 2.7100 0.3200 2.8000 0.6850 ;
        RECT 3.2300 0.3200 3.3200 0.6850 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9000 0.3500 1.2500 ;
        RECT 0.2500 0.8000 0.5650 0.9000 ;
        RECT 0.4650 0.5800 0.5650 0.8000 ;
        RECT 0.4650 0.4800 0.9750 0.5800 ;
        RECT 0.8750 0.5800 0.9750 1.1600 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END G

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2550 0.5500 1.3950 ;
        RECT 0.4500 1.0450 0.5850 1.2550 ;
    END
    ANTENNAGATEAREA 0.0747 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4450 1.4500 3.1500 1.5500 ;
        RECT 2.4450 1.5500 2.5450 1.8800 ;
        RECT 2.9650 1.5500 3.0650 1.8800 ;
        RECT 3.0500 0.9500 3.1500 1.4500 ;
        RECT 2.4500 0.8500 3.1500 0.9500 ;
        RECT 2.4500 0.5200 2.5400 0.8500 ;
        RECT 2.9650 0.5200 3.0650 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.3350 1.9400 0.4350 2.0800 ;
        RECT 1.6800 1.7700 1.7700 2.0800 ;
        RECT 2.1900 1.7700 2.2800 2.0800 ;
        RECT 2.7100 1.7700 2.8000 2.0800 ;
        RECT 3.2300 1.7700 3.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6750 0.6800 0.7650 1.6150 ;
      RECT 0.0700 1.7300 0.9500 1.8200 ;
      RECT 0.8600 1.3800 0.9500 1.7300 ;
      RECT 0.8600 1.2900 1.2550 1.3800 ;
      RECT 1.1650 0.8200 1.2550 1.2900 ;
      RECT 0.0700 1.8200 0.1700 1.9350 ;
      RECT 0.0700 0.6950 0.1600 1.7300 ;
      RECT 0.0700 0.4850 0.2100 0.6950 ;
      RECT 1.3650 0.9450 1.8750 1.0350 ;
      RECT 1.7850 1.0350 1.8750 1.2000 ;
      RECT 1.0600 1.5700 1.1500 1.9100 ;
      RECT 1.0600 1.4800 1.4550 1.5700 ;
      RECT 1.3650 1.0350 1.4550 1.4800 ;
      RECT 1.3650 0.7100 1.4550 0.9450 ;
      RECT 1.0650 0.6200 1.4550 0.7100 ;
      RECT 2.0550 1.0900 2.8000 1.1800 ;
      RECT 1.5450 1.1550 1.6350 1.3200 ;
      RECT 1.9400 1.4100 2.0300 1.7500 ;
      RECT 1.5450 1.3200 2.1450 1.4100 ;
      RECT 2.0550 1.1800 2.1450 1.3200 ;
      RECT 2.0550 0.8550 2.1450 1.0900 ;
      RECT 1.9400 0.7650 2.1450 0.8550 ;
      RECT 1.9400 0.4450 2.0300 0.7650 ;
  END
END LATQN_X4M_A12TH

MACRO LATQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 1.6000 0.3200 1.7000 0.7400 ;
        RECT 1.9650 0.3200 2.0650 0.7750 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9000 0.5750 1.2500 ;
    END
    ANTENNAGATEAREA 0.0291 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2300 0.6050 2.3500 1.7200 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9150 0.3500 1.4500 ;
        RECT 0.2500 1.4500 0.5500 1.5500 ;
        RECT 0.4500 1.5500 0.5500 1.8200 ;
        RECT 0.4500 1.8200 1.2500 1.9200 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.9700 1.5350 2.0600 2.0800 ;
        RECT 1.4600 1.5300 1.5500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6650 1.5650 0.8400 1.6550 ;
      RECT 0.6650 0.7700 0.7550 1.5650 ;
      RECT 0.6650 0.6800 0.8850 0.7700 ;
      RECT 0.2050 0.4800 1.0650 0.5700 ;
      RECT 0.9750 0.5700 1.0650 0.8900 ;
      RECT 0.8450 0.8900 1.3200 0.9800 ;
      RECT 0.8450 0.9800 0.9350 1.4550 ;
      RECT 0.0500 1.7100 0.2400 1.8000 ;
      RECT 0.0500 0.7550 0.1400 1.7100 ;
      RECT 0.0500 0.6650 0.2950 0.7550 ;
      RECT 0.2050 0.5700 0.2950 0.6650 ;
      RECT 1.0500 1.1100 1.9500 1.2000 ;
      RECT 1.4100 0.7600 1.5000 1.1100 ;
      RECT 1.1550 0.6700 1.5000 0.7600 ;
      RECT 0.9350 1.5900 1.1400 1.6800 ;
      RECT 1.0500 1.2000 1.1400 1.5900 ;
      RECT 1.1550 0.5450 1.2450 0.6700 ;
      RECT 1.3500 1.3200 2.1350 1.4100 ;
      RECT 2.0450 0.9550 2.1350 1.3200 ;
      RECT 1.5900 0.8650 2.1350 0.9550 ;
  END
END LATQ_X0P5M_A12TH

MACRO LATQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.4450 ;
        RECT 0.6650 0.3200 0.8350 0.5400 ;
        RECT 1.9000 0.3200 2.0000 0.6450 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5150 0.1700 1.7200 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7700 1.2100 1.9500 1.4600 ;
        RECT 1.7700 1.0500 1.8750 1.2100 ;
    END
    ANTENNAGATEAREA 0.0675 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9500 2.1550 1.2800 ;
        RECT 1.7100 0.8500 2.1550 0.9500 ;
        RECT 1.7100 0.5800 1.8100 0.8500 ;
        RECT 1.3450 0.4800 1.8100 0.5800 ;
        RECT 1.3450 0.5800 1.4350 1.2400 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3400 1.7650 0.4300 2.0800 ;
        RECT 0.7050 1.7400 0.7950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6150 1.3200 0.8400 1.4100 ;
      RECT 0.7500 0.9200 0.8400 1.3200 ;
      RECT 0.6150 0.8300 0.8400 0.9200 ;
      RECT 1.1550 1.6650 1.2450 1.9150 ;
      RECT 0.9300 1.5750 1.2450 1.6650 ;
      RECT 0.9300 0.7200 1.0200 1.5750 ;
      RECT 0.3450 0.6300 1.2550 0.7200 ;
      RECT 1.1650 0.4300 1.2550 0.6300 ;
      RECT 0.3450 0.7200 0.4350 1.2300 ;
      RECT 1.5250 0.6950 1.6150 1.7200 ;
      RECT 1.3450 1.8300 2.1400 1.9200 ;
      RECT 2.0500 1.7550 2.1400 1.8300 ;
      RECT 2.0500 1.6650 2.3550 1.7550 ;
      RECT 2.2650 0.5600 2.3550 1.6650 ;
      RECT 2.1650 0.4700 2.3550 0.5600 ;
      RECT 1.1100 0.8400 1.2000 1.3550 ;
      RECT 1.3450 1.4450 1.4350 1.8300 ;
      RECT 1.1100 1.3550 1.4350 1.4450 ;
  END
END LATQ_X1M_A12TH

MACRO LATQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.3350 0.3200 0.5200 0.5400 ;
        RECT 0.8350 0.3200 1.0450 0.3700 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 0.8300 0.8500 0.9500 ;
        RECT 0.7500 0.9500 0.8500 1.3400 ;
        RECT 0.5550 1.3400 0.8500 1.4400 ;
    END
    ANTENNADIFFAREA 0.3432 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.1050 2.1500 1.5500 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9800 2.3500 1.1900 ;
        RECT 2.0500 0.8800 2.3500 0.9800 ;
        RECT 2.0500 0.5700 2.1500 0.8800 ;
        RECT 1.6500 0.4800 2.1500 0.5700 ;
        RECT 1.6500 0.5700 1.7400 0.8500 ;
        RECT 1.5700 0.8500 1.7400 0.9400 ;
        RECT 1.5700 0.9400 1.6600 1.2400 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 2.0700 2.0350 2.2400 2.0800 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8950 1.7700 0.9850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6300 1.0800 0.7200 ;
      RECT 0.9900 0.7200 1.0800 1.2000 ;
      RECT 0.0800 0.7200 0.1700 1.4700 ;
      RECT 1.4900 1.6500 1.5800 1.9700 ;
      RECT 0.2800 1.5600 1.5800 1.6500 ;
      RECT 1.1700 0.7500 1.2600 1.5600 ;
      RECT 1.1700 0.6600 1.5200 0.7500 ;
      RECT 1.4300 0.5300 1.5200 0.6600 ;
      RECT 0.2800 1.1700 0.3700 1.5600 ;
      RECT 0.2800 1.0800 0.6500 1.1700 ;
      RECT 1.8500 0.6650 1.9400 1.7100 ;
      RECT 1.6700 1.8200 2.5400 1.9100 ;
      RECT 2.4000 1.3050 2.5400 1.8200 ;
      RECT 2.4500 0.7900 2.5400 1.3050 ;
      RECT 2.4000 0.5800 2.5400 0.7900 ;
      RECT 1.3700 0.8400 1.4600 1.3700 ;
      RECT 1.6700 1.4600 1.7600 1.8200 ;
      RECT 1.3700 1.3700 1.7600 1.4600 ;
  END
END LATQ_X2M_A12TH

MACRO LATQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6850 ;
        RECT 0.8600 0.3200 0.9500 0.4650 ;
        RECT 1.2150 0.3200 1.4250 0.5400 ;
        RECT 2.5050 0.3200 2.6050 0.4200 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4450 1.0200 2.5500 1.4550 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9000 2.7750 1.1900 ;
        RECT 2.4500 0.8000 2.7750 0.9000 ;
        RECT 2.4500 0.6100 2.5500 0.8000 ;
        RECT 2.0400 0.5100 2.5500 0.6100 ;
        RECT 2.0400 0.6100 2.1400 1.1050 ;
        RECT 1.9200 1.1050 2.1400 1.2050 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END G

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4500 0.6900 1.5500 ;
        RECT 0.0800 1.5500 0.1700 1.8800 ;
        RECT 0.6000 1.5500 0.6900 1.8800 ;
        RECT 0.2500 0.9500 0.3500 1.4500 ;
        RECT 0.0800 0.8500 0.6900 0.9500 ;
        RECT 0.0800 0.5200 0.1700 0.8500 ;
        RECT 0.6000 0.5200 0.6900 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 2.5100 1.8400 2.6000 2.0800 ;
        RECT 0.3400 1.7700 0.4300 2.0800 ;
        RECT 0.8600 1.7700 0.9500 2.0800 ;
        RECT 1.2750 1.5200 1.3650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1400 1.3200 1.3700 1.4100 ;
      RECT 1.2800 0.9400 1.3700 1.3200 ;
      RECT 1.1400 0.8500 1.3700 0.9400 ;
      RECT 1.8700 1.6300 1.9600 1.9600 ;
      RECT 1.4600 1.5400 1.9600 1.6300 ;
      RECT 0.9000 0.6300 1.9200 0.7200 ;
      RECT 1.8300 0.4300 1.9200 0.6300 ;
      RECT 1.4600 0.7200 1.5500 1.5400 ;
      RECT 0.9000 0.7200 0.9900 1.0800 ;
      RECT 0.4700 1.0800 0.9900 1.1700 ;
      RECT 2.2500 0.7050 2.3400 1.5000 ;
      RECT 2.0500 1.6600 2.9550 1.7500 ;
      RECT 2.8100 1.3000 2.9550 1.6600 ;
      RECT 2.8650 0.6150 2.9550 1.3000 ;
      RECT 2.8050 0.4250 2.9550 0.6150 ;
      RECT 1.6900 0.8100 1.7800 1.3400 ;
      RECT 2.0500 1.4300 2.1400 1.6600 ;
      RECT 1.6900 1.3400 2.1400 1.4300 ;
  END
END LATQ_X3M_A12TH

MACRO LATRPQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 1.0150 0.3200 1.1050 0.4350 ;
        RECT 2.2250 0.3200 2.3750 0.9000 ;
        RECT 0.9350 0.4350 1.1050 0.5250 ;
        RECT 1.0150 0.5250 1.1050 0.9250 ;
    END
  END VSS

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7250 0.5550 0.9500 ;
        RECT 0.4500 0.9500 0.6000 1.1850 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.2300 2.3500 1.6650 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1950 1.9500 1.3900 ;
        RECT 1.6950 1.0100 1.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.4250 0.1700 1.8450 ;
        RECT 0.0450 0.5200 0.1500 1.4250 ;
        RECT 0.0450 0.4300 0.2400 0.5200 ;
    END
    ANTENNADIFFAREA 0.1377 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.0450 1.7550 1.1350 2.0800 ;
        RECT 0.3500 1.6350 0.4400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8150 1.5050 1.1800 1.5650 ;
      RECT 0.2650 1.4750 1.1800 1.5050 ;
      RECT 0.8150 1.5650 0.9050 1.8950 ;
      RECT 0.2650 1.4150 0.9050 1.4750 ;
      RECT 0.6900 0.5150 0.7800 1.4150 ;
      RECT 0.6150 0.4250 0.8250 0.5150 ;
      RECT 0.2650 1.0450 0.3550 1.4150 ;
      RECT 1.2700 0.7600 1.7050 0.8500 ;
      RECT 1.2700 1.8150 1.6350 1.9050 ;
      RECT 1.2700 1.2850 1.3600 1.8150 ;
      RECT 0.8700 1.1950 1.3600 1.2850 ;
      RECT 1.2700 0.8500 1.3600 1.1950 ;
      RECT 1.9250 1.6500 2.1300 1.7400 ;
      RECT 2.0400 0.8650 2.1300 1.6500 ;
      RECT 1.8150 0.7750 2.1300 0.8650 ;
      RECT 1.7250 1.8300 2.7500 1.9200 ;
      RECT 2.6600 0.8600 2.7500 1.8300 ;
      RECT 2.5500 0.7700 2.7500 0.8600 ;
      RECT 1.4500 0.9600 1.5400 1.5400 ;
      RECT 1.7250 1.6300 1.8150 1.8300 ;
      RECT 1.4500 1.5400 1.8150 1.6300 ;
  END
END LATRPQN_X0P5M_A12TH

MACRO LATRPQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 1.0050 0.3200 1.0950 0.9300 ;
        RECT 2.2200 0.3200 2.3900 0.8850 ;
    END
  END VSS

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7250 0.5500 0.9500 ;
        RECT 0.4500 0.9500 0.6000 1.1850 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.1900 2.3500 1.6100 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6750 1.0600 1.9500 1.2300 ;
        RECT 1.8500 0.8100 1.9500 1.0600 ;
    END
    ANTENNAGATEAREA 0.0594 ;
  END G

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4250 0.1700 1.8450 ;
        RECT 0.0500 0.8950 0.1500 1.4250 ;
        RECT 0.0500 0.4800 0.1700 0.8950 ;
    END
    ANTENNADIFFAREA 0.27625 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.2350 2.0100 2.4450 2.0800 ;
        RECT 0.3100 1.8950 0.4800 2.0800 ;
        RECT 1.0450 1.6900 1.1350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8150 1.5450 1.1800 1.5650 ;
      RECT 0.2650 1.4750 1.1800 1.5450 ;
      RECT 0.8150 1.5650 0.9050 1.9050 ;
      RECT 0.2650 1.4550 0.9050 1.4750 ;
      RECT 0.6900 0.5150 0.7800 1.4550 ;
      RECT 0.6150 0.4250 0.8250 0.5150 ;
      RECT 0.2650 1.0450 0.3550 1.4550 ;
      RECT 1.2700 0.6750 1.7600 0.7650 ;
      RECT 1.2700 1.7500 1.6350 1.8400 ;
      RECT 1.2700 1.2850 1.3600 1.7500 ;
      RECT 0.8700 1.1950 1.3600 1.2850 ;
      RECT 1.2700 0.7650 1.3600 1.1950 ;
      RECT 1.9250 1.6450 2.1300 1.7350 ;
      RECT 2.0400 0.6900 2.1300 1.6450 ;
      RECT 1.8700 0.6000 2.1300 0.6900 ;
      RECT 1.7250 1.8300 2.7500 1.9200 ;
      RECT 2.6600 0.8400 2.7500 1.8300 ;
      RECT 2.5500 0.7500 2.7500 0.8400 ;
      RECT 1.4500 0.9400 1.5400 1.4300 ;
      RECT 1.7250 1.5200 1.8150 1.8300 ;
      RECT 1.4500 1.4300 1.8150 1.5200 ;
  END
END LATRPQN_X1M_A12TH

MACRO INV_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.1550 0.3200 0.2550 0.8250 ;
        RECT 0.6400 0.3200 0.8100 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.4150 1.2500 1.1500 1.3500 ;
        RECT 0.4150 0.8500 1.1500 0.9500 ;
        RECT 0.4150 1.3500 0.5150 1.7350 ;
        RECT 0.9350 1.3500 1.0350 1.7350 ;
        RECT 0.4150 0.4400 0.5150 0.8500 ;
        RECT 0.9350 0.4400 1.0350 0.8500 ;
    END
    ANTENNADIFFAREA 0.552825 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.1550 1.7700 0.2550 2.0800 ;
        RECT 0.6750 1.7700 0.7750 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3100 1.0500 0.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.2457 ;
  END A
END INV_X3B_A12TH

MACRO INV_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6350 ;
        RECT 0.6100 0.3200 0.7100 0.6350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9500 0.9700 1.2500 ;
        RECT 0.3500 1.2500 0.9700 1.3500 ;
        RECT 0.3500 0.8500 0.9700 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7200 ;
        RECT 0.8700 1.3500 0.9700 1.7200 ;
        RECT 0.3500 0.4900 0.4500 0.8500 ;
        RECT 0.8700 0.4900 0.9700 0.8500 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.0500 0.7300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2925 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
    END
  END VDD
END INV_X3M_A12TH

MACRO INV_X3P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1550 0.3200 0.2550 0.8050 ;
        RECT 0.6400 0.3200 0.8100 0.7100 ;
        RECT 1.1600 0.3200 1.3300 0.7100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4200 1.0500 1.0300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2868 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1550 1.6550 0.2550 2.0800 ;
        RECT 0.6750 1.6550 0.7750 2.0800 ;
        RECT 1.1950 1.6550 1.2950 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.2500 ;
        RECT 0.4150 1.2500 1.3500 1.3500 ;
        RECT 0.4150 0.8500 1.3500 0.9500 ;
        RECT 0.4150 1.3500 0.5150 1.7200 ;
        RECT 0.9350 1.3500 1.0350 1.7200 ;
        RECT 0.4150 0.4450 0.5150 0.8500 ;
        RECT 0.9350 0.4450 1.0350 0.8500 ;
    END
    ANTENNADIFFAREA 0.478 ;
  END Y
END INV_X3P5B_A12TH

MACRO INV_X3P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1000 0.3200 0.2000 0.7250 ;
        RECT 0.6200 0.3200 0.7200 0.7250 ;
        RECT 1.1400 0.3200 1.2400 0.7250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1000 1.6550 0.2000 2.0800 ;
        RECT 0.6200 1.6550 0.7200 2.0800 ;
        RECT 1.1400 1.6550 1.2400 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.0500 0.8450 1.1500 ;
    END
    ANTENNAGATEAREA 0.3408 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.3600 1.2500 1.1500 1.3500 ;
        RECT 0.3600 0.8500 1.1500 0.9500 ;
        RECT 0.3600 1.3500 0.4600 1.7200 ;
        RECT 0.8800 1.3500 0.9800 1.7200 ;
        RECT 0.3600 0.4850 0.4600 0.8500 ;
        RECT 0.8800 0.4850 0.9800 0.8500 ;
    END
    ANTENNADIFFAREA 0.568 ;
  END Y
END INV_X3P5M_A12TH

MACRO INV_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.7200 ;
        RECT 0.6450 0.3200 0.7350 0.7100 ;
        RECT 1.1600 0.3200 1.2600 0.7100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.3276 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 1.4500 1.1500 1.5500 ;
        RECT 0.3800 1.5500 0.4800 1.8800 ;
        RECT 0.9000 1.5500 1.0000 1.8800 ;
        RECT 1.0500 0.9500 1.1500 1.4500 ;
        RECT 0.3800 0.8500 1.1500 0.9500 ;
        RECT 0.3800 0.4400 0.4800 0.8500 ;
        RECT 0.9000 0.4400 1.0000 0.8500 ;
    END
    ANTENNADIFFAREA 0.546 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1200 2.0600 0.7400 2.0800 ;
        RECT 1.1600 1.7500 1.2600 2.0800 ;
        RECT 0.1200 1.7500 0.2200 2.0600 ;
        RECT 0.6400 1.7500 0.7400 2.0600 ;
    END
  END VDD
END INV_X4B_A12TH

MACRO INV_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6350 ;
        RECT 0.6100 0.3200 0.7100 0.6350 ;
        RECT 1.1300 0.3200 1.2300 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 0.7500 1.1500 ;
    END
    ANTENNAGATEAREA 0.39 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.3500 1.2500 1.1500 1.3500 ;
        RECT 0.3500 0.8500 1.1500 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7200 ;
        RECT 0.8700 1.3500 0.9700 1.7250 ;
        RECT 0.3500 0.4900 0.4500 0.8500 ;
        RECT 0.8700 0.4900 0.9700 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y
END INV_X4M_A12TH

MACRO INV_X5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.1000 0.3200 0.2000 0.8250 ;
        RECT 0.5850 0.3200 0.7550 0.7300 ;
        RECT 1.1050 0.3200 1.2750 0.7300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.2500 ;
        RECT 0.3600 1.2500 1.5500 1.3500 ;
        RECT 0.3600 0.8500 1.5500 0.9500 ;
        RECT 0.3600 1.3500 0.4600 1.7350 ;
        RECT 0.8800 1.3500 0.9800 1.7350 ;
        RECT 1.4000 1.3500 1.5500 1.7350 ;
        RECT 0.3600 0.4400 0.4600 0.8500 ;
        RECT 0.8800 0.4400 0.9800 0.8500 ;
        RECT 1.4050 0.4400 1.5500 0.8500 ;
    END
    ANTENNADIFFAREA 0.7917 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.1000 1.7700 0.2000 2.0800 ;
        RECT 0.6200 1.7700 0.7200 2.0800 ;
        RECT 1.1400 1.7700 1.2400 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.0500 1.2200 1.1500 ;
    END
    ANTENNAGATEAREA 0.4095 ;
  END A
END INV_X5B_A12TH

MACRO INV_X5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.1050 0.3200 0.2050 0.6350 ;
        RECT 0.6300 0.3200 0.7300 0.6350 ;
        RECT 1.1500 0.3200 1.2500 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.1050 1.7700 0.2050 2.0800 ;
        RECT 0.6300 1.7700 0.7300 2.0800 ;
        RECT 1.1500 1.7700 1.2500 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.3700 1.2500 1.5100 1.3500 ;
        RECT 0.3700 0.8500 1.5100 0.9500 ;
        RECT 0.3700 1.3500 0.4700 1.7200 ;
        RECT 0.8900 1.3500 0.9900 1.7200 ;
        RECT 1.4100 1.3500 1.5100 1.7200 ;
        RECT 0.3700 0.4900 0.4700 0.8500 ;
        RECT 0.8900 0.4900 0.9900 0.8500 ;
        RECT 1.4100 0.4900 1.5100 0.8500 ;
    END
    ANTENNADIFFAREA 0.934375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 1.0500 0.8250 1.1500 ;
    END
    ANTENNAGATEAREA 0.4875 ;
  END A
END INV_X5M_A12TH

MACRO INV_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1750 0.3200 0.2750 0.8250 ;
        RECT 0.6600 0.3200 0.8300 0.7100 ;
        RECT 1.1800 0.3200 1.3500 0.7100 ;
        RECT 1.7000 0.3200 1.8700 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.2500 ;
        RECT 0.4350 1.2500 1.7500 1.3500 ;
        RECT 0.4350 0.8500 1.7500 0.9500 ;
        RECT 0.4350 1.3500 0.5350 1.7200 ;
        RECT 0.9550 1.3500 1.0550 1.7200 ;
        RECT 1.4750 1.3500 1.5750 1.7200 ;
        RECT 1.4750 0.4550 1.5750 0.8500 ;
        RECT 0.4350 0.4400 0.5350 0.8500 ;
        RECT 0.9550 0.4400 1.0550 0.8500 ;
    END
    ANTENNADIFFAREA 0.819 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1750 1.7700 0.2750 2.0800 ;
        RECT 0.6950 1.7700 0.7950 2.0800 ;
        RECT 1.2150 1.7700 1.3150 2.0800 ;
        RECT 1.7350 1.7700 1.8350 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3350 1.0500 1.1450 1.1500 ;
    END
    ANTENNAGATEAREA 0.4914 ;
  END A
END INV_X6B_A12TH

MACRO INV_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1250 0.3200 0.2250 0.6350 ;
        RECT 0.6450 0.3200 0.7450 0.6350 ;
        RECT 1.1650 0.3200 1.2650 0.6350 ;
        RECT 1.6850 0.3200 1.7850 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5000 1.0500 1.3000 1.1500 ;
    END
    ANTENNAGATEAREA 0.585 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.1250 1.7700 0.2250 2.0800 ;
        RECT 0.6450 1.7700 0.7450 2.0800 ;
        RECT 1.1650 1.7700 1.2650 2.0800 ;
        RECT 1.6800 1.7700 1.7900 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4250 1.3500 1.5500 1.7200 ;
        RECT 0.3850 1.2500 1.5500 1.3500 ;
        RECT 0.3850 1.3500 0.4850 1.7200 ;
        RECT 0.9050 1.3500 1.0050 1.7200 ;
        RECT 1.4500 0.9500 1.5500 1.2500 ;
        RECT 0.3850 0.8500 1.5500 0.9500 ;
        RECT 0.3850 0.4900 0.4850 0.8500 ;
        RECT 0.9050 0.4900 1.0050 0.8500 ;
        RECT 1.4250 0.4900 1.5500 0.8500 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y
END INV_X6M_A12TH

MACRO INV_X7P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.1100 1.7150 0.2100 2.0800 ;
        RECT 0.6300 1.7150 0.7300 2.0800 ;
        RECT 1.1500 1.7150 1.2500 2.0800 ;
        RECT 1.6700 1.7150 1.7700 2.0800 ;
        RECT 2.1900 1.7150 2.2900 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1100 0.3200 0.2100 0.8200 ;
        RECT 0.5950 0.3200 0.7650 0.7000 ;
        RECT 1.1150 0.3200 1.2850 0.7000 ;
        RECT 1.6350 0.3200 1.8050 0.7000 ;
        RECT 2.1550 0.3200 2.3250 0.7000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0450 0.9550 2.1550 1.2450 ;
        RECT 0.3700 1.2450 2.1550 1.3550 ;
        RECT 0.3700 0.8450 2.1550 0.9550 ;
        RECT 0.3700 1.3550 0.4700 1.7200 ;
        RECT 0.8900 1.3550 0.9900 1.7200 ;
        RECT 1.4050 1.3550 1.5150 1.7200 ;
        RECT 1.9300 1.3550 2.0300 1.7200 ;
        RECT 0.3700 0.4400 0.4700 0.8450 ;
        RECT 0.8900 0.4400 0.9900 0.8450 ;
        RECT 1.4100 0.4400 1.5100 0.8450 ;
        RECT 1.9300 0.4400 2.0300 0.8450 ;
    END
    ANTENNADIFFAREA 1.028 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.0500 1.6300 1.1500 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END A
END INV_X7P5B_A12TH

MACRO INV_X7P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.6550 ;
        RECT 0.6000 0.3200 0.7000 0.6750 ;
        RECT 1.1200 0.3200 1.2200 0.6750 ;
        RECT 1.6400 0.3200 1.7400 0.6750 ;
        RECT 2.1600 0.3200 2.2600 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.0800 1.7150 0.1800 2.0800 ;
        RECT 0.6000 1.7150 0.7000 2.0800 ;
        RECT 1.1200 1.7150 1.2200 2.0800 ;
        RECT 1.6400 1.7150 1.7400 2.0800 ;
        RECT 2.1600 1.7150 2.2600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6400 0.9200 1.7600 1.4400 ;
        RECT 0.3400 1.4400 2.0000 1.5600 ;
        RECT 0.3400 0.8000 2.0000 0.9200 ;
        RECT 0.3400 1.5600 0.4400 1.8700 ;
        RECT 0.8600 1.5600 0.9600 1.8700 ;
        RECT 1.3800 1.5600 1.4800 1.8700 ;
        RECT 1.9000 1.5600 2.0000 1.8700 ;
        RECT 0.3400 0.4900 0.4400 0.8000 ;
        RECT 0.8600 0.4900 0.9600 0.8000 ;
        RECT 1.3800 0.4900 1.4800 0.8000 ;
        RECT 1.9000 0.4900 2.0000 0.8000 ;
    END
    ANTENNADIFFAREA 1.224 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 1.0500 1.3400 1.1500 ;
    END
    ANTENNAGATEAREA 0.7344 ;
  END A
END INV_X7P5M_A12TH

MACRO INV_X9B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8050 ;
        RECT 0.5600 0.3200 0.7300 0.6800 ;
        RECT 1.0800 0.3200 1.2500 0.6800 ;
        RECT 1.6000 0.3200 1.7700 0.6800 ;
        RECT 2.1200 0.3200 2.2900 0.6800 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 1.0500 1.8250 1.1500 ;
    END
    ANTENNAGATEAREA 0.7371 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 0.5950 1.7700 0.6950 2.0800 ;
        RECT 1.1150 1.7700 1.2150 2.0800 ;
        RECT 1.6350 1.7700 1.7350 2.0800 ;
        RECT 2.1550 1.7700 2.2550 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3350 1.4350 2.5150 1.5650 ;
        RECT 0.3350 1.5650 0.4350 1.8650 ;
        RECT 0.8550 1.5650 0.9550 1.8650 ;
        RECT 1.3750 1.5650 1.4750 1.8650 ;
        RECT 1.8950 1.5650 1.9950 1.8650 ;
        RECT 2.4150 1.5650 2.5150 1.8650 ;
        RECT 2.3850 0.9300 2.5150 1.4350 ;
        RECT 0.3350 0.8000 2.5150 0.9300 ;
        RECT 0.3350 0.4400 0.4350 0.8000 ;
        RECT 0.8550 0.4400 0.9550 0.8000 ;
        RECT 1.3750 0.4400 1.4750 0.8000 ;
        RECT 1.8950 0.4400 1.9950 0.8000 ;
        RECT 2.4150 0.4400 2.5150 0.8000 ;
    END
    ANTENNADIFFAREA 1.3104 ;
  END Y
END INV_X9B_A12TH

MACRO INV_X9M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.6350 ;
        RECT 0.6000 0.3200 0.7000 0.6350 ;
        RECT 1.1200 0.3200 1.2200 0.6350 ;
        RECT 1.6400 0.3200 1.7400 0.6350 ;
        RECT 2.1600 0.3200 2.2600 0.6350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6350 0.9200 1.7650 1.4350 ;
        RECT 0.3400 1.4350 2.5200 1.5650 ;
        RECT 0.3400 0.7900 2.5200 0.9200 ;
        RECT 0.3400 1.5650 0.4400 1.8650 ;
        RECT 0.8600 1.5650 0.9600 1.8650 ;
        RECT 1.3800 1.5650 1.4800 1.8650 ;
        RECT 1.9000 1.5650 2.0000 1.8650 ;
        RECT 2.4200 1.5650 2.5200 1.8650 ;
        RECT 0.3400 0.4900 0.4400 0.7900 ;
        RECT 0.8600 0.4900 0.9600 0.7900 ;
        RECT 1.3800 0.4900 1.4800 0.7900 ;
        RECT 1.9000 0.4900 2.0000 0.7900 ;
        RECT 2.4200 0.4900 2.5200 0.7900 ;
    END
    ANTENNADIFFAREA 1.568125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5100 1.0500 1.3450 1.1500 ;
    END
    ANTENNAGATEAREA 0.8775 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.0800 1.7700 0.1800 2.0800 ;
        RECT 0.6000 1.7700 0.7000 2.0800 ;
        RECT 1.1200 1.7700 1.2200 2.0800 ;
        RECT 1.6400 1.7700 1.7400 2.0800 ;
        RECT 2.1600 1.7700 2.2600 2.0800 ;
    END
  END VDD
END INV_X9M_A12TH

MACRO LATNQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 1.6500 0.3200 1.7600 0.8000 ;
        RECT 2.1650 0.3200 2.2650 0.9600 ;
    END
  END VSS

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.4950 0.5500 1.8300 ;
        RECT 0.4500 1.8300 1.1250 1.9200 ;
        RECT 0.2700 1.3850 0.5500 1.4950 ;
        RECT 0.2700 1.0700 0.3700 1.3850 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END GN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5900 0.9000 0.7500 1.2750 ;
    END
    ANTENNAGATEAREA 0.0291 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4250 1.3950 2.5500 1.7200 ;
        RECT 2.4250 0.5500 2.5250 1.3950 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 1.6650 1.6000 1.7650 2.0800 ;
        RECT 2.1650 1.3200 2.2650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7300 1.6150 0.9300 1.7100 ;
      RECT 0.8400 0.7800 0.9300 1.6150 ;
      RECT 0.7100 0.6800 0.9300 0.7800 ;
      RECT 1.2450 1.2650 1.3350 1.4900 ;
      RECT 1.0200 1.1750 1.3350 1.2650 ;
      RECT 1.0200 0.5700 1.1100 1.1750 ;
      RECT 0.0800 0.4800 1.1100 0.5700 ;
      RECT 0.0800 0.5700 0.1700 1.7950 ;
      RECT 1.4250 0.8900 1.8350 0.9800 ;
      RECT 1.7450 0.9800 1.8350 1.0800 ;
      RECT 1.1400 1.6200 1.5150 1.7100 ;
      RECT 1.4250 0.9800 1.5150 1.6200 ;
      RECT 1.4250 0.7800 1.5150 0.8900 ;
      RECT 1.2000 0.6900 1.5150 0.7800 ;
      RECT 1.2000 0.5900 1.3000 0.6900 ;
      RECT 1.9400 1.0900 2.2500 1.1950 ;
      RECT 1.6050 1.4000 1.7000 1.4900 ;
      RECT 1.6050 1.3050 2.0350 1.4000 ;
      RECT 1.9350 1.4000 2.0350 1.7850 ;
      RECT 1.9400 1.1950 2.0350 1.3050 ;
      RECT 1.9400 0.6050 2.0350 1.0900 ;
  END
END LATNQN_X0P5M_A12TH

MACRO LATNQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 1.6500 0.3200 1.7600 0.7800 ;
        RECT 2.1650 0.3200 2.2650 0.6550 ;
    END
  END VSS

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.4850 0.5500 1.8300 ;
        RECT 0.4500 1.8300 1.1200 1.9200 ;
        RECT 0.2700 1.3750 0.5500 1.4850 ;
        RECT 0.2700 0.9950 0.3700 1.3750 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END GN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5900 0.8950 0.7500 1.2650 ;
    END
    ANTENNAGATEAREA 0.0372 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4250 1.3950 2.5500 1.8550 ;
        RECT 2.4250 0.4900 2.5250 1.3950 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 2.1650 1.7650 2.2650 2.0800 ;
        RECT 1.6550 1.6000 1.7550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7250 1.6150 0.9300 1.7100 ;
      RECT 0.8400 0.7800 0.9300 1.6150 ;
      RECT 0.7200 0.6800 0.9300 0.7800 ;
      RECT 1.2250 1.2650 1.3150 1.5100 ;
      RECT 1.0200 1.1750 1.3150 1.2650 ;
      RECT 1.0200 0.5700 1.1100 1.1750 ;
      RECT 0.0800 0.4800 1.1100 0.5700 ;
      RECT 0.0800 0.5700 0.1700 1.7950 ;
      RECT 1.4050 0.8700 1.8250 0.9600 ;
      RECT 1.7350 0.9600 1.8250 1.0600 ;
      RECT 1.1300 1.6350 1.4950 1.7250 ;
      RECT 1.4050 0.9600 1.4950 1.6350 ;
      RECT 1.4050 0.7800 1.4950 0.8700 ;
      RECT 1.2000 0.6900 1.4950 0.7800 ;
      RECT 1.2000 0.5900 1.3000 0.6900 ;
      RECT 1.9200 1.0900 2.2500 1.1950 ;
      RECT 1.5850 1.4000 1.6800 1.4900 ;
      RECT 1.5850 1.3050 2.0150 1.4000 ;
      RECT 1.9150 1.4000 2.0150 1.9800 ;
      RECT 1.9200 1.1950 2.0150 1.3050 ;
      RECT 1.9200 0.6050 2.0150 1.0900 ;
  END
END LATNQN_X1M_A12TH

MACRO LATNQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.9200 0.3200 1.0100 0.4400 ;
        RECT 0.3350 0.3200 0.4400 0.5300 ;
        RECT 2.0600 0.3200 2.2600 0.3900 ;
        RECT 0.8000 0.4400 1.0100 0.5300 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9700 1.0100 2.1500 1.2350 ;
        RECT 1.9700 0.8650 2.0700 1.0100 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.2950 1.6800 1.3950 ;
        RECT 1.5900 1.3950 1.6800 1.8300 ;
        RECT 1.2500 0.8000 1.3500 1.2950 ;
        RECT 1.5900 1.8300 2.3400 1.9200 ;
        RECT 2.2500 1.0300 2.3400 1.8300 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9800 0.9500 1.4450 ;
        RECT 0.5950 1.4450 0.9500 1.5450 ;
        RECT 0.5900 0.8800 0.9500 0.9800 ;
        RECT 0.5950 1.5450 0.6950 1.8650 ;
        RECT 0.5900 0.8000 0.7000 0.8800 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.8500 1.7750 0.9600 2.0800 ;
        RECT 0.3350 1.4650 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4850 1.1050 0.6850 1.2050 ;
      RECT 0.0550 1.2650 0.5750 1.3550 ;
      RECT 0.4850 1.2050 0.5750 1.2650 ;
      RECT 0.0550 1.3550 0.1750 1.7400 ;
      RECT 0.0550 0.6150 0.1450 1.2650 ;
      RECT 0.0550 0.4100 0.1700 0.6150 ;
      RECT 1.4100 1.6500 1.5000 1.7850 ;
      RECT 1.0400 1.5600 1.5000 1.6500 ;
      RECT 0.2600 0.6200 1.4500 0.7100 ;
      RECT 1.3600 0.4300 1.4500 0.6200 ;
      RECT 1.0400 0.7100 1.1300 1.5600 ;
      RECT 0.2600 0.7100 0.3500 1.1750 ;
      RECT 1.7900 0.7600 1.8800 1.7400 ;
      RECT 1.7400 0.6600 1.9350 0.7600 ;
      RECT 1.5400 0.4800 2.5200 0.5700 ;
      RECT 2.4300 0.5700 2.5200 1.8700 ;
      RECT 1.5400 0.5700 1.6300 0.9600 ;
  END
END LATNQN_X2M_A12TH

MACRO LATNQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.2750 0.3200 0.4900 0.4200 ;
        RECT 0.8000 0.3200 1.0100 0.4200 ;
        RECT 1.3250 0.3200 1.4950 0.5300 ;
        RECT 2.5600 0.3200 2.6600 0.6050 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3700 1.2000 2.5500 1.3950 ;
        RECT 2.3700 1.0150 2.4650 1.2000 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.3000 2.1000 1.3900 ;
        RECT 1.6500 0.9700 1.7500 1.3000 ;
        RECT 2.0100 1.3900 2.1000 1.8300 ;
        RECT 1.6500 0.8000 1.8100 0.9700 ;
        RECT 2.0100 1.8300 2.7400 1.9200 ;
        RECT 2.6500 1.0300 2.7400 1.8300 ;
    END
    ANTENNAGATEAREA 0.0786 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5950 1.4500 1.2150 1.5500 ;
        RECT 0.5950 1.5500 0.6950 1.8950 ;
        RECT 1.1150 1.5500 1.2150 1.8950 ;
        RECT 1.1150 0.9300 1.2150 1.4500 ;
        RECT 0.5400 0.8300 1.2900 0.9300 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 2.4150 2.0750 2.5850 2.0800 ;
        RECT 0.8500 1.7750 0.9600 2.0800 ;
        RECT 1.3450 1.7000 1.4450 2.0800 ;
        RECT 0.3350 1.6250 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4850 1.1050 0.9100 1.2050 ;
      RECT 0.0550 1.3600 0.1750 1.7400 ;
      RECT 0.0550 0.8150 0.1450 1.2700 ;
      RECT 0.0550 0.4100 0.1700 0.8150 ;
      RECT 0.0550 1.2700 0.5750 1.3600 ;
      RECT 0.4850 1.2050 0.5750 1.2700 ;
      RECT 1.8300 1.5900 1.9200 1.9100 ;
      RECT 1.4400 1.5000 1.9200 1.5900 ;
      RECT 0.2600 0.6200 1.9050 0.7100 ;
      RECT 1.8150 0.4300 1.9050 0.6200 ;
      RECT 1.4400 0.7100 1.5300 1.5000 ;
      RECT 0.2600 0.7100 0.3550 1.1800 ;
      RECT 2.1900 0.7100 2.2800 1.7200 ;
      RECT 2.8300 0.8350 2.9200 1.9350 ;
      RECT 2.3800 0.7450 2.9200 0.8350 ;
      RECT 2.8300 0.4100 2.9200 0.7450 ;
      RECT 2.3800 0.5700 2.4700 0.7450 ;
      RECT 1.9950 0.4800 2.4700 0.5700 ;
      RECT 1.9950 0.5700 2.0850 1.0650 ;
  END
END LATNQN_X3M_A12TH

MACRO LATNQN_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.2750 0.3200 0.4900 0.4200 ;
        RECT 0.8000 0.3200 1.0100 0.4200 ;
        RECT 1.4150 0.3200 1.5850 0.5300 ;
        RECT 2.7600 0.3200 2.8600 0.6050 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5700 1.2000 2.7500 1.3950 ;
        RECT 2.5700 1.0150 2.6650 1.2000 ;
    END
    ANTENNAGATEAREA 0.0747 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.2800 2.3000 1.3900 ;
        RECT 2.2100 1.3900 2.3000 1.8300 ;
        RECT 1.8500 0.9700 1.9500 1.2800 ;
        RECT 2.2100 1.8300 2.9400 1.9200 ;
        RECT 1.8500 0.8000 1.9900 0.9700 ;
        RECT 2.8500 1.0150 2.9400 1.8300 ;
    END
    ANTENNAGATEAREA 0.0948 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5950 1.4500 1.2150 1.5500 ;
        RECT 0.5950 1.5500 0.6950 1.8950 ;
        RECT 1.1150 1.5500 1.2150 1.8950 ;
        RECT 1.1150 0.9200 1.2150 1.4500 ;
        RECT 0.5400 0.8200 1.2750 0.9200 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.8500 1.7750 0.9600 2.0800 ;
        RECT 0.3350 1.7700 0.4350 2.0800 ;
        RECT 1.3750 1.7700 1.4750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4850 1.1050 0.9100 1.2050 ;
      RECT 0.0550 1.3600 0.1750 1.7400 ;
      RECT 0.0550 0.8150 0.1450 1.2700 ;
      RECT 0.0550 0.4100 0.1700 0.8150 ;
      RECT 0.0550 1.2700 0.5750 1.3600 ;
      RECT 0.4850 1.2050 0.5750 1.2700 ;
      RECT 2.0300 1.5900 2.1200 1.9100 ;
      RECT 1.6400 1.5000 2.1200 1.5900 ;
      RECT 0.2600 0.6200 2.0850 0.7100 ;
      RECT 1.9950 0.4100 2.0850 0.6200 ;
      RECT 1.6400 0.7100 1.7300 1.5000 ;
      RECT 0.2600 0.7100 0.3550 1.1800 ;
      RECT 2.3900 0.7100 2.4800 1.7200 ;
      RECT 3.0300 0.8350 3.1200 1.9350 ;
      RECT 2.5800 0.7450 3.1200 0.8350 ;
      RECT 3.0300 0.4100 3.1200 0.7450 ;
      RECT 2.5800 0.5700 2.6700 0.7450 ;
      RECT 2.1950 0.4800 2.6700 0.5700 ;
      RECT 2.1950 0.5700 2.2850 1.1700 ;
  END
END LATNQN_X4M_A12TH

MACRO LATNQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3600 0.3200 0.4500 0.4900 ;
        RECT 0.6200 0.3200 0.7900 0.5250 ;
        RECT 1.9150 0.3200 2.0050 0.6300 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 0.9500 1.9550 1.2250 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0450 0.8100 1.1550 1.3500 ;
        RECT 1.0450 1.3500 1.4500 1.4600 ;
        RECT 1.3400 1.4600 1.4500 1.8200 ;
        RECT 1.3400 1.8200 1.9500 1.9200 ;
        RECT 1.8500 1.7100 1.9500 1.8200 ;
        RECT 1.8500 1.6100 2.1400 1.7100 ;
        RECT 2.0400 1.2550 2.1400 1.6100 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5250 0.1700 1.7200 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.9000 2.0100 1.9900 2.0800 ;
        RECT 0.3600 1.8750 0.4500 2.0800 ;
        RECT 0.5900 1.8750 0.7600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6600 1.2200 0.7500 1.4650 ;
      RECT 0.6600 1.0500 0.8100 1.2200 ;
      RECT 0.6600 0.8000 0.7500 1.0500 ;
      RECT 0.4600 1.6450 1.2300 1.7350 ;
      RECT 1.1400 1.5650 1.2300 1.6450 ;
      RECT 0.4600 0.6200 1.2100 0.7100 ;
      RECT 1.1200 0.4100 1.2100 0.6200 ;
      RECT 0.4600 1.2050 0.5500 1.6450 ;
      RECT 0.2600 1.0350 0.5500 1.2050 ;
      RECT 0.4600 0.7100 0.5500 1.0350 ;
      RECT 1.5400 0.6900 1.6300 1.7100 ;
      RECT 1.7350 0.7700 2.3200 0.8600 ;
      RECT 2.2300 0.8600 2.3200 1.7650 ;
      RECT 2.2300 0.4100 2.3200 0.7700 ;
      RECT 1.3450 0.4800 1.8250 0.5700 ;
      RECT 1.7350 0.5700 1.8250 0.7700 ;
      RECT 1.2650 1.1300 1.4350 1.2200 ;
      RECT 1.3450 0.5700 1.4350 1.1300 ;
  END
END LATNQ_X0P5M_A12TH

MACRO LATNQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.4150 ;
        RECT 0.5450 0.3200 0.7150 0.5250 ;
        RECT 1.9350 0.3200 2.0250 0.6000 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 0.9500 1.9500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0675 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.6100 2.1400 1.7100 ;
        RECT 1.6500 1.7100 1.7500 1.8200 ;
        RECT 2.0400 1.2550 2.1400 1.6100 ;
        RECT 1.2900 1.8200 1.7500 1.9200 ;
        RECT 1.2900 1.4000 1.3800 1.8200 ;
        RECT 1.1350 1.3100 1.3800 1.4000 ;
        RECT 1.1350 0.8100 1.2250 1.3100 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.4900 0.1700 1.7200 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.8600 1.8550 1.9500 2.0800 ;
        RECT 0.5350 1.7800 0.6250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6500 1.3500 0.7400 1.4700 ;
      RECT 0.6500 1.2600 0.8450 1.3500 ;
      RECT 0.7550 0.8900 0.8450 1.2600 ;
      RECT 0.5900 0.8000 0.8450 0.8900 ;
      RECT 1.1100 1.5800 1.2000 1.9650 ;
      RECT 0.9350 1.4900 1.2000 1.5800 ;
      RECT 0.2650 0.6200 1.2100 0.7100 ;
      RECT 1.1200 0.4100 1.2100 0.6200 ;
      RECT 0.9350 0.7100 1.0250 1.4900 ;
      RECT 0.2650 1.0200 0.5550 1.1900 ;
      RECT 0.2650 0.7100 0.3550 1.0200 ;
      RECT 1.4700 1.4100 1.7050 1.5000 ;
      RECT 1.6150 1.0400 1.7050 1.4100 ;
      RECT 1.5550 0.9500 1.7050 1.0400 ;
      RECT 1.4700 1.5000 1.5600 1.7100 ;
      RECT 1.5550 0.6900 1.6450 0.9500 ;
      RECT 1.7350 0.7700 2.3200 0.8600 ;
      RECT 2.2300 0.8600 2.3200 1.7550 ;
      RECT 2.2300 0.4100 2.3200 0.7700 ;
      RECT 1.3350 1.1300 1.5050 1.2200 ;
      RECT 1.3350 0.5700 1.4250 1.1300 ;
      RECT 1.3350 0.4800 1.8250 0.5700 ;
      RECT 1.7350 0.5700 1.8250 0.7700 ;
  END
END LATNQ_X1M_A12TH

MACRO LATNQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3600 0.3200 0.5300 0.5200 ;
        RECT 0.9200 0.3200 1.0900 0.5200 ;
        RECT 2.3100 0.3200 2.4000 0.3950 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9000 0.7500 1.5000 ;
        RECT 0.6000 0.7900 0.8100 0.9000 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7350 2.3650 1.1100 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.2500 1.9500 1.3500 ;
        RECT 1.8600 1.3500 1.9500 1.6500 ;
        RECT 1.4500 1.1400 1.5400 1.2500 ;
        RECT 1.8600 1.6500 2.4500 1.7500 ;
        RECT 2.3500 1.4400 2.4500 1.6500 ;
        RECT 2.3500 1.3400 2.5650 1.4400 ;
        RECT 2.4650 1.1300 2.5650 1.3400 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END GN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.2900 1.8450 2.5000 2.0800 ;
        RECT 0.4000 1.7900 0.4900 2.0800 ;
        RECT 0.9350 1.7900 1.0250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6100 1.1600 0.7000 ;
      RECT 1.0700 0.7000 1.1600 1.1950 ;
      RECT 0.0800 0.7000 0.1700 1.4700 ;
      RECT 1.6800 1.7000 1.7700 1.9900 ;
      RECT 0.4700 1.6100 1.7700 1.7000 ;
      RECT 1.2500 0.9600 1.7600 1.0500 ;
      RECT 1.6700 0.4300 1.7600 0.9600 ;
      RECT 1.2500 1.0500 1.3400 1.6100 ;
      RECT 0.4700 1.2100 0.5600 1.6100 ;
      RECT 0.2600 1.0400 0.5600 1.2100 ;
      RECT 2.0500 1.3800 2.2400 1.5000 ;
      RECT 2.0500 0.6650 2.1400 1.3800 ;
      RECT 2.6300 1.6550 2.7200 1.9800 ;
      RECT 2.6300 1.5750 2.7450 1.6550 ;
      RECT 2.6550 0.7500 2.7450 1.5750 ;
      RECT 2.6300 0.5750 2.7450 0.7500 ;
      RECT 1.8500 0.4850 2.7450 0.5750 ;
      RECT 1.8500 0.5750 1.9400 1.1000 ;
  END
END LATNQ_X2M_A12TH

MACRO LATNQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6850 ;
        RECT 0.8600 0.3200 0.9500 0.4650 ;
        RECT 1.1750 0.3200 1.2650 0.5200 ;
        RECT 2.4300 0.3200 2.5200 0.4350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3650 0.8500 2.6000 0.9500 ;
        RECT 2.3650 0.9500 2.4650 1.1400 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3600 1.2800 2.7500 1.3900 ;
        RECT 2.3600 1.3900 2.4600 1.6500 ;
        RECT 2.6500 1.0600 2.7500 1.2800 ;
        RECT 1.9700 1.6500 2.4600 1.7500 ;
        RECT 1.9700 1.2300 2.0700 1.6500 ;
        RECT 1.5400 1.1200 2.0700 1.2300 ;
        RECT 1.5400 0.9200 1.6300 1.1200 ;
    END
    ANTENNAGATEAREA 0.0894 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 0.6950 1.5500 ;
        RECT 0.0750 1.5500 0.1750 1.8600 ;
        RECT 0.5950 1.5500 0.6950 1.8600 ;
        RECT 0.0750 0.9900 0.1750 1.4500 ;
        RECT 0.0750 0.8900 0.6950 0.9900 ;
        RECT 0.0750 0.5400 0.1750 0.8900 ;
        RECT 0.5950 0.5400 0.6950 0.8900 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 1.2250 1.9700 1.3150 2.0800 ;
        RECT 0.3400 1.7700 0.4300 2.0800 ;
        RECT 0.8600 1.7700 0.9500 2.0800 ;
        RECT 2.5700 1.4800 2.6600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1800 1.6400 1.2900 1.8800 ;
      RECT 1.1800 1.5500 1.4350 1.6400 ;
      RECT 1.1800 1.0000 1.2700 1.5500 ;
      RECT 1.1600 0.8100 1.2700 1.0000 ;
      RECT 1.7900 1.4600 1.8800 1.9100 ;
      RECT 1.3600 1.3700 1.8800 1.4600 ;
      RECT 1.3600 0.7000 1.8800 0.7800 ;
      RECT 0.8450 0.6900 1.8800 0.7000 ;
      RECT 1.7900 0.4100 1.8800 0.6900 ;
      RECT 1.3600 0.7800 1.4500 1.3700 ;
      RECT 0.8450 0.6100 1.4500 0.6900 ;
      RECT 0.8450 0.7000 0.9350 1.0800 ;
      RECT 0.3250 1.0800 0.9350 1.1700 ;
      RECT 2.1700 0.7050 2.2600 1.5000 ;
      RECT 2.8300 1.4400 2.9450 1.8300 ;
      RECT 2.8550 0.7000 2.9450 1.4400 ;
      RECT 2.3700 0.6150 2.9450 0.7000 ;
      RECT 1.9700 0.6100 2.9450 0.6150 ;
      RECT 1.9700 0.6150 2.0600 0.9200 ;
      RECT 1.8100 0.9200 2.0600 1.0100 ;
      RECT 1.9700 0.5250 2.4600 0.6100 ;
  END
END LATNQ_X3M_A12TH

MACRO LATNRPQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.9350 0.3200 1.0250 0.5750 ;
        RECT 0.3400 0.3200 0.4300 0.7550 ;
        RECT 2.3300 0.3200 2.5000 0.6900 ;
        RECT 0.9350 0.5750 1.1300 0.6750 ;
        RECT 1.0400 0.6750 1.1300 0.7800 ;
    END
  END VSS

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9100 0.6000 1.1900 ;
    END
    ANTENNAGATEAREA 0.0309 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1300 1.0500 2.5500 1.1500 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8700 1.5500 1.3850 ;
        RECT 1.4500 1.3850 1.8300 1.4750 ;
        RECT 1.7400 1.4750 1.8300 1.8300 ;
        RECT 1.7400 1.8300 2.2300 1.9200 ;
        RECT 2.1400 1.5900 2.2300 1.8300 ;
        RECT 2.1400 1.5000 2.5300 1.5900 ;
        RECT 2.4400 1.3400 2.5300 1.5000 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END GN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.5150 0.1700 0.7350 ;
        RECT 0.0500 0.7350 0.1500 1.7200 ;
        RECT 0.0500 1.7200 0.1700 1.9900 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.3400 1.7950 0.4300 2.0800 ;
        RECT 2.3200 1.7150 2.4100 2.0800 ;
        RECT 1.0400 1.5700 1.1300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2450 1.3800 1.1600 1.4700 ;
      RECT 1.0700 1.2900 1.1600 1.3800 ;
      RECT 0.2450 1.2650 0.3350 1.3800 ;
      RECT 0.8150 1.4700 0.9050 1.9900 ;
      RECT 0.6900 0.5050 0.7800 1.3800 ;
      RECT 0.6150 0.4150 0.8250 0.5050 ;
      RECT 1.5600 1.6750 1.6500 1.7900 ;
      RECT 1.2500 1.5850 1.6500 1.6750 ;
      RECT 1.2500 0.6900 1.5900 0.7800 ;
      RECT 1.5000 0.5900 1.5900 0.6900 ;
      RECT 1.2500 1.0950 1.3400 1.5850 ;
      RECT 0.8700 1.0050 1.3400 1.0950 ;
      RECT 1.2500 0.7800 1.3400 1.0050 ;
      RECT 0.8700 0.8850 0.9600 1.0050 ;
      RECT 1.9400 0.7700 2.0300 1.7400 ;
      RECT 1.8600 0.6800 2.0300 0.7700 ;
      RECT 2.6300 1.6600 2.7400 1.8800 ;
      RECT 2.6500 0.8700 2.7400 1.6600 ;
      RECT 2.1200 0.7800 2.7400 0.8700 ;
      RECT 2.6300 0.5550 2.7400 0.7800 ;
      RECT 2.1200 0.5700 2.2100 0.7800 ;
      RECT 1.6800 0.4800 2.2100 0.5700 ;
      RECT 1.6800 0.5700 1.7700 1.2800 ;
  END
END LATNRPQN_X0P5M_A12TH

MACRO LATNRPQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.9750 0.3200 2.4500 0.3250 ;
        RECT 0.3200 0.3200 0.5300 0.5300 ;
        RECT 0.9750 0.3250 1.0750 0.8250 ;
        RECT 2.2400 0.3250 2.4500 0.4350 ;
    END
  END VSS

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 1.6500 2.5400 1.7500 ;
        RECT 1.7950 1.2400 1.8850 1.6500 ;
        RECT 2.4500 1.0050 2.5400 1.6500 ;
        RECT 1.3850 1.1500 1.8850 1.2400 ;
        RECT 1.3850 1.0300 1.4750 1.1500 ;
    END
    ANTENNAGATEAREA 0.0609 ;
  END GN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1550 0.9850 2.3500 1.2050 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3300 0.8500 0.6000 0.9500 ;
        RECT 0.5100 0.6800 0.6000 0.8500 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END R

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9200 0.1500 1.2900 ;
        RECT 0.0500 1.2900 0.1750 1.7000 ;
        RECT 0.0500 0.5150 0.1750 0.9200 ;
    END
    ANTENNADIFFAREA 0.263575 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.2700 1.8700 2.4400 2.0800 ;
        RECT 0.9950 1.7450 1.2000 2.0800 ;
        RECT 0.3450 1.6850 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8050 1.5100 1.2550 1.6350 ;
      RECT 0.8050 1.2650 0.8950 1.5100 ;
      RECT 0.3400 1.1750 0.8950 1.2650 ;
      RECT 0.7100 0.5400 0.8000 1.1750 ;
      RECT 0.6400 0.4500 0.8500 0.5400 ;
      RECT 0.3400 1.1500 0.4300 1.1750 ;
      RECT 0.2400 1.0600 0.4300 1.1500 ;
      RECT 1.6150 1.4200 1.7050 1.8050 ;
      RECT 1.1850 1.3300 1.7050 1.4200 ;
      RECT 1.1850 0.8300 1.6300 0.9200 ;
      RECT 1.5400 0.6250 1.6300 0.8300 ;
      RECT 1.1850 1.0650 1.2750 1.3300 ;
      RECT 0.8900 0.9750 1.2750 1.0650 ;
      RECT 1.1850 0.9200 1.2750 0.9750 ;
      RECT 1.9750 0.8000 2.0650 1.5400 ;
      RECT 1.9200 0.7100 2.1100 0.8000 ;
      RECT 1.7200 0.5300 2.7200 0.6200 ;
      RECT 2.6300 0.6200 2.7200 1.5550 ;
      RECT 1.7200 0.6200 1.8100 1.0400 ;
  END
END LATNRPQN_X1M_A12TH

MACRO LATNRPQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.1400 0.3200 0.2300 0.7900 ;
        RECT 0.7500 0.3200 0.8400 0.5600 ;
        RECT 1.2700 0.3200 1.3600 0.6200 ;
        RECT 2.5350 0.3200 2.6250 0.8050 ;
    END
  END VSS

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8700 1.7700 1.2500 ;
        RECT 1.6500 1.2500 2.0850 1.3500 ;
        RECT 1.9950 1.3500 2.0850 1.8300 ;
        RECT 1.9950 1.8300 2.5500 1.9200 ;
        RECT 2.4600 1.7900 2.5500 1.8300 ;
        RECT 2.4600 1.7000 2.7400 1.7900 ;
        RECT 2.6500 1.1550 2.7400 1.7000 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END GN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5850 0.8400 0.7900 0.9500 ;
        RECT 0.5850 0.9500 0.7050 1.1150 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3750 1.1900 2.5500 1.4000 ;
        RECT 2.4500 1.4000 2.5500 1.5900 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9300 1.1500 1.4250 ;
        RECT 0.9000 1.4250 1.1500 1.5150 ;
        RECT 1.0100 0.8400 1.1500 0.9300 ;
        RECT 1.0100 0.5600 1.1000 0.8400 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 2.5100 2.0100 2.6000 2.0800 ;
        RECT 1.2750 1.8350 1.3650 2.0800 ;
        RECT 0.6400 1.8200 0.7300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4050 1.2250 0.9450 1.3150 ;
      RECT 0.8550 1.0200 0.9450 1.2250 ;
      RECT 0.0450 0.9700 0.1350 1.5850 ;
      RECT 0.1200 1.6750 0.2100 1.9550 ;
      RECT 0.0450 1.5850 0.2100 1.6750 ;
      RECT 0.0450 0.8800 0.4950 0.9700 ;
      RECT 0.4050 0.9700 0.4950 1.2250 ;
      RECT 0.4050 0.4450 0.4950 0.8800 ;
      RECT 1.8150 1.7150 1.9050 1.8350 ;
      RECT 0.5650 1.6250 1.9050 1.7150 ;
      RECT 1.4500 0.6100 1.9050 0.7000 ;
      RECT 1.8150 0.4300 1.9050 0.6100 ;
      RECT 1.4500 0.7000 1.5400 1.6250 ;
      RECT 0.5650 1.4950 0.6550 1.6250 ;
      RECT 0.2250 1.4050 0.6550 1.4950 ;
      RECT 0.2250 1.0800 0.3150 1.4050 ;
      RECT 2.1750 1.6300 2.3600 1.7200 ;
      RECT 2.1750 0.6800 2.2650 1.6300 ;
      RECT 2.8300 1.0050 2.9200 1.9750 ;
      RECT 2.3550 0.9150 2.9200 1.0050 ;
      RECT 2.8300 0.5800 2.9200 0.9150 ;
      RECT 1.9950 0.5700 2.0850 1.1300 ;
      RECT 2.3550 0.5700 2.4450 0.9150 ;
      RECT 1.9950 0.4800 2.4450 0.5700 ;
  END
END LATNRPQN_X2M_A12TH

MACRO INV_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.1300 0.3200 0.2300 0.8550 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9750 0.3500 1.3950 ;
    END
    ANTENNAGATEAREA 0.0411 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8700 0.5500 1.5000 ;
        RECT 0.4100 1.5000 0.5500 1.6000 ;
        RECT 0.4150 0.6600 0.5500 0.8700 ;
        RECT 0.4100 1.6000 0.5100 1.9100 ;
    END
    ANTENNADIFFAREA 0.119875 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.1300 1.5450 0.2300 2.0800 ;
    END
  END VDD
END INV_X0P5B_A12TH

MACRO INV_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.1300 0.3200 0.2300 0.8550 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9800 0.3500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8700 0.5500 1.5000 ;
        RECT 0.4100 1.5000 0.5500 1.6000 ;
        RECT 0.4100 0.7700 0.5500 0.8700 ;
        RECT 0.4100 1.6000 0.5100 1.9100 ;
        RECT 0.4100 0.4600 0.5100 0.7700 ;
    END
    ANTENNADIFFAREA 0.142625 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.1300 1.5450 0.2300 2.0800 ;
    END
  END VDD
END INV_X0P5M_A12TH

MACRO INV_X0P6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.7750 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7800 0.5500 1.5000 ;
        RECT 0.3550 1.5000 0.5500 1.6000 ;
        RECT 0.3000 0.6800 0.5500 0.7800 ;
        RECT 0.3550 1.6000 0.4550 1.9300 ;
    END
    ANTENNADIFFAREA 0.16605 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9150 0.3500 1.3350 ;
    END
    ANTENNAGATEAREA 0.0486 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0950 1.5200 0.1950 2.0800 ;
    END
  END VDD
END INV_X0P6B_A12TH

MACRO INV_X0P6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.8800 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8750 0.5500 1.5250 ;
        RECT 0.3550 1.5250 0.5500 1.6250 ;
        RECT 0.3550 0.7750 0.5500 0.8750 ;
        RECT 0.3550 1.6250 0.4550 1.9600 ;
        RECT 0.3550 0.4400 0.4550 0.7750 ;
    END
    ANTENNADIFFAREA 0.168875 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9850 0.3500 1.4050 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0950 1.5300 0.1950 2.0800 ;
    END
  END VDD
END INV_X0P6M_A12TH

MACRO INV_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.6300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.6900 0.5500 1.3850 ;
        RECT 0.3550 1.3850 0.5500 1.4850 ;
        RECT 0.3000 0.5900 0.5500 0.6900 ;
        RECT 0.3550 1.4850 0.4550 1.8250 ;
    END
    ANTENNADIFFAREA 0.19885 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8250 0.3500 1.2450 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0950 1.5300 0.1950 2.0800 ;
    END
  END VDD
END INV_X0P7B_A12TH

MACRO INV_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1800 0.8350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8750 0.5500 1.5200 ;
        RECT 0.3550 1.5200 0.5500 1.6200 ;
        RECT 0.3550 0.7750 0.5500 0.8750 ;
        RECT 0.3550 1.6200 0.4550 1.9600 ;
        RECT 0.3550 0.4400 0.4550 0.7750 ;
    END
    ANTENNADIFFAREA 0.202125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9850 0.3500 1.4050 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0950 1.5300 0.1950 2.0800 ;
    END
  END VDD
END INV_X0P7M_A12TH

MACRO INV_X0P8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8750 0.5500 1.5400 ;
        RECT 0.3500 1.5400 0.5500 1.6400 ;
        RECT 0.3550 0.7750 0.5500 0.8750 ;
        RECT 0.3500 1.6400 0.4500 1.9600 ;
        RECT 0.3550 0.4450 0.4550 0.7750 ;
    END
    ANTENNADIFFAREA 0.23575 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0000 0.3500 1.4200 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0750 1.6800 0.1750 2.0800 ;
    END
  END VDD
END INV_X0P8B_A12TH

MACRO INV_X0P8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7450 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8800 0.5500 1.5350 ;
        RECT 0.3500 1.5350 0.5500 1.6350 ;
        RECT 0.3550 0.7800 0.5500 0.8800 ;
        RECT 0.3500 1.6350 0.4500 1.9600 ;
        RECT 0.3550 0.4400 0.4550 0.7800 ;
    END
    ANTENNADIFFAREA 0.238875 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0000 0.3500 1.4250 ;
    END
    ANTENNAGATEAREA 0.0819 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0750 1.6500 0.1750 2.0800 ;
    END
  END VDD
END INV_X0P8M_A12TH

MACRO INV_X11B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.7750 ;
        RECT 0.6050 0.3200 0.7750 0.6500 ;
        RECT 1.1250 0.3200 1.2950 0.6500 ;
        RECT 1.6450 0.3200 1.8150 0.6500 ;
        RECT 2.1650 0.3200 2.3350 0.6500 ;
        RECT 2.6850 0.3200 2.8550 0.6500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 1.4200 3.0750 1.5800 ;
        RECT 0.3800 1.5800 0.4800 1.8500 ;
        RECT 0.9000 1.5800 1.0000 1.8500 ;
        RECT 1.4200 1.5800 1.5200 1.8500 ;
        RECT 1.9400 1.5800 2.0400 1.8500 ;
        RECT 2.4600 1.5800 2.5600 1.8500 ;
        RECT 2.9850 1.5800 3.0750 1.8500 ;
        RECT 2.8200 0.9300 2.9800 1.4200 ;
        RECT 0.3850 0.7700 3.0750 0.9300 ;
        RECT 0.3850 0.4400 0.4750 0.7700 ;
        RECT 0.9050 0.4400 0.9950 0.7700 ;
        RECT 1.4250 0.4400 1.5150 0.7700 ;
        RECT 1.9450 0.4400 2.0350 0.7700 ;
        RECT 2.4650 0.4400 2.5550 0.7700 ;
        RECT 2.9850 0.4400 3.0750 0.7700 ;
    END
    ANTENNADIFFAREA 1.6107 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.1200 1.7700 0.2200 2.0800 ;
        RECT 0.6400 1.7700 0.7400 2.0800 ;
        RECT 1.1600 1.7700 1.2600 2.0800 ;
        RECT 1.6800 1.7700 1.7800 2.0800 ;
        RECT 2.2000 1.7700 2.3000 2.0800 ;
        RECT 2.7200 1.7700 2.8200 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 2.1750 1.1500 ;
    END
    ANTENNAGATEAREA 0.9009 ;
  END A
END INV_X11B_A12TH

MACRO INV_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1000 0.3200 0.2000 0.6350 ;
        RECT 0.6200 0.3200 0.7200 0.6350 ;
        RECT 1.1400 0.3200 1.2400 0.6350 ;
        RECT 1.6600 0.3200 1.7600 0.6350 ;
        RECT 2.1800 0.3200 2.2800 0.6350 ;
        RECT 2.7000 0.3200 2.8000 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 1.0500 1.9000 1.1600 ;
    END
    ANTENNAGATEAREA 1.0725 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2200 0.9200 2.3800 1.4200 ;
        RECT 0.3600 1.4200 3.0600 1.5800 ;
        RECT 0.3600 0.7600 3.0600 0.9200 ;
        RECT 0.3600 1.5800 0.4600 1.8500 ;
        RECT 0.8800 1.5800 0.9800 1.8500 ;
        RECT 1.4000 1.5800 1.5000 1.8500 ;
        RECT 1.9200 1.5800 2.0200 1.8500 ;
        RECT 2.4400 1.5800 2.5400 1.8500 ;
        RECT 2.9600 1.5800 3.0600 1.8500 ;
        RECT 0.3600 0.4900 0.4600 0.7600 ;
        RECT 0.8800 0.4900 0.9800 0.7600 ;
        RECT 1.4000 0.4900 1.5000 0.7600 ;
        RECT 1.9200 0.4900 2.0200 0.7600 ;
        RECT 2.4400 0.4900 2.5400 0.7600 ;
        RECT 2.9600 0.4900 3.0600 0.7600 ;
    END
    ANTENNADIFFAREA 1.909375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.1000 1.7700 0.2000 2.0800 ;
        RECT 0.6200 1.7700 0.7200 2.0800 ;
        RECT 1.1400 1.7700 1.2400 2.0800 ;
        RECT 1.6600 1.7700 1.7600 2.0800 ;
        RECT 2.1800 1.7700 2.2800 2.0800 ;
        RECT 2.7000 1.7700 2.8000 2.0800 ;
    END
  END VDD
END INV_X11M_A12TH

MACRO INV_X13B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.1600 0.3200 0.2600 0.7850 ;
        RECT 0.6450 0.3200 0.8150 0.6600 ;
        RECT 1.1650 0.3200 1.3350 0.6600 ;
        RECT 1.6850 0.3200 1.8550 0.6600 ;
        RECT 2.2050 0.3200 2.3750 0.6600 ;
        RECT 2.7250 0.3200 2.8950 0.6600 ;
        RECT 3.2450 0.3200 3.4150 0.6600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4200 1.4100 3.6400 1.5900 ;
        RECT 0.4200 1.5900 0.5200 1.8400 ;
        RECT 0.9400 1.5900 1.0400 1.8400 ;
        RECT 1.4600 1.5900 1.5600 1.8400 ;
        RECT 1.9800 1.5900 2.0800 1.8400 ;
        RECT 2.5000 1.5900 2.6000 1.8400 ;
        RECT 3.0200 1.5900 3.1200 1.8400 ;
        RECT 3.5400 1.5900 3.6400 1.8400 ;
        RECT 3.2100 0.9300 3.3900 1.4100 ;
        RECT 0.4200 0.7500 3.6350 0.9300 ;
        RECT 0.4200 0.4400 0.5200 0.7500 ;
        RECT 0.9400 0.4400 1.0400 0.7500 ;
        RECT 1.4600 0.4400 1.5600 0.7500 ;
        RECT 1.9800 0.4400 2.0800 0.7500 ;
        RECT 2.5000 0.4400 2.6000 0.7500 ;
        RECT 3.0200 0.4400 3.1200 0.7500 ;
        RECT 3.5450 0.4400 3.6350 0.7500 ;
    END
    ANTENNADIFFAREA 1.917825 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.1600 1.7700 0.2600 2.0800 ;
        RECT 0.6800 1.7700 0.7800 2.0800 ;
        RECT 1.2000 1.7700 1.3000 2.0800 ;
        RECT 1.7200 1.7700 1.8200 2.0800 ;
        RECT 2.2400 1.7700 2.3400 2.0800 ;
        RECT 2.7600 1.7700 2.8600 2.0800 ;
        RECT 3.2800 1.7700 3.3800 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5900 1.0500 2.7500 1.1500 ;
    END
    ANTENNAGATEAREA 1.0647 ;
  END A
END INV_X13B_A12TH

MACRO INV_X13M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.1450 0.3200 0.2450 0.6150 ;
        RECT 0.6650 0.3200 0.7650 0.6150 ;
        RECT 1.1850 0.3200 1.2850 0.6150 ;
        RECT 1.7050 0.3200 1.8050 0.6150 ;
        RECT 2.2250 0.3200 2.3250 0.6150 ;
        RECT 2.7450 0.3200 2.8450 0.6150 ;
        RECT 3.2650 0.3200 3.3650 0.6150 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.0500 2.4550 1.1500 ;
    END
    ANTENNAGATEAREA 1.2675 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.1450 1.7700 0.2450 2.0800 ;
        RECT 0.6650 1.7700 0.7650 2.0800 ;
        RECT 1.1850 1.7700 1.2850 2.0800 ;
        RECT 1.7050 1.7700 1.8050 2.0800 ;
        RECT 2.2250 1.7700 2.3250 2.0800 ;
        RECT 2.7450 1.7700 2.8450 2.0800 ;
        RECT 3.2650 1.7700 3.3650 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8100 0.9200 2.9900 1.4100 ;
        RECT 0.4050 1.4100 3.6250 1.5900 ;
        RECT 0.4050 0.7400 3.6250 0.9200 ;
        RECT 0.4050 1.5900 0.5050 1.8400 ;
        RECT 0.9250 1.5900 1.0250 1.8400 ;
        RECT 1.4450 1.5900 1.5450 1.8400 ;
        RECT 1.9650 1.5900 2.0650 1.8400 ;
        RECT 2.4850 1.5900 2.5850 1.8400 ;
        RECT 3.0050 1.5900 3.1050 1.8400 ;
        RECT 3.5250 1.5900 3.6250 1.8400 ;
        RECT 0.4050 0.4900 0.5050 0.7400 ;
        RECT 0.9250 0.4900 1.0250 0.7400 ;
        RECT 1.4450 0.4900 1.5450 0.7400 ;
        RECT 1.9650 0.4900 2.0650 0.7400 ;
        RECT 2.4850 0.4900 2.5850 0.7400 ;
        RECT 3.0050 0.4900 3.1050 0.7400 ;
        RECT 3.5250 0.4900 3.6250 0.7400 ;
    END
    ANTENNADIFFAREA 2.234375 ;
  END Y
END INV_X13M_A12TH

MACRO INV_X16B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1700 0.3200 0.2700 0.7550 ;
        RECT 0.6550 0.3200 0.8250 0.6300 ;
        RECT 1.1750 0.3200 1.3450 0.6300 ;
        RECT 1.6950 0.3200 1.8650 0.6300 ;
        RECT 2.2150 0.3200 2.3850 0.6300 ;
        RECT 2.7350 0.3200 2.9050 0.6300 ;
        RECT 3.2550 0.3200 3.4250 0.6300 ;
        RECT 3.7750 0.3200 3.9450 0.6300 ;
        RECT 4.3350 0.3200 4.4250 0.7550 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9900 0.9400 4.2100 1.3900 ;
        RECT 0.4350 1.3900 4.2100 1.6100 ;
        RECT 0.4300 0.7200 4.2100 0.9400 ;
        RECT 0.4350 1.6100 0.5250 1.8200 ;
        RECT 0.9550 1.6100 1.0450 1.8200 ;
        RECT 1.4750 1.6100 1.5650 1.8200 ;
        RECT 1.9950 1.6100 2.0850 1.8200 ;
        RECT 2.5150 1.6100 2.6050 1.8200 ;
        RECT 3.0350 1.6100 3.1250 1.8200 ;
        RECT 3.5550 1.6100 3.6450 1.8200 ;
        RECT 4.0700 1.6100 4.2100 1.8200 ;
        RECT 0.4300 0.4200 0.5300 0.7200 ;
        RECT 0.9500 0.4200 1.0500 0.7200 ;
        RECT 1.4700 0.4200 1.5700 0.7200 ;
        RECT 1.9900 0.4200 2.0900 0.7200 ;
        RECT 2.5100 0.4200 2.6100 0.7200 ;
        RECT 3.0300 0.4200 3.1300 0.7200 ;
        RECT 3.5500 0.4200 3.6500 0.7200 ;
        RECT 4.0700 0.4200 4.2100 0.7200 ;
    END
    ANTENNADIFFAREA 2.184 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1700 1.7700 0.2700 2.0800 ;
        RECT 0.6900 1.7700 0.7900 2.0800 ;
        RECT 1.2100 1.7700 1.3100 2.0800 ;
        RECT 1.7300 1.7700 1.8300 2.0800 ;
        RECT 2.2500 1.7700 2.3500 2.0800 ;
        RECT 2.7700 1.7700 2.8700 2.0800 ;
        RECT 3.2900 1.7700 3.3900 2.0800 ;
        RECT 3.8100 1.7700 3.9100 2.0800 ;
        RECT 4.3300 1.7700 4.4300 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 3.3400 1.1500 ;
    END
    ANTENNAGATEAREA 1.3104 ;
  END A
END INV_X16B_A12TH

MACRO INV_X16M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1700 0.3200 0.2700 0.6100 ;
        RECT 0.6900 0.3200 0.7900 0.5900 ;
        RECT 1.2100 0.3200 1.3100 0.5900 ;
        RECT 1.7300 0.3200 1.8300 0.5900 ;
        RECT 2.2500 0.3200 2.3500 0.5900 ;
        RECT 2.7700 0.3200 2.8700 0.5900 ;
        RECT 3.2900 0.3200 3.3900 0.5900 ;
        RECT 3.8100 0.3200 3.9100 0.5900 ;
        RECT 4.3300 0.3200 4.4300 0.6100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5900 0.9300 3.8100 1.3900 ;
        RECT 0.4200 1.3900 4.1800 1.6100 ;
        RECT 0.4200 0.7100 4.1800 0.9300 ;
        RECT 0.4200 1.6100 0.5400 1.8200 ;
        RECT 0.9400 1.6100 1.0600 1.8200 ;
        RECT 1.4600 1.6100 1.5800 1.8200 ;
        RECT 1.9800 1.6100 2.1000 1.8200 ;
        RECT 2.5000 1.6100 2.6200 1.8200 ;
        RECT 3.0200 1.6100 3.1400 1.8200 ;
        RECT 3.5400 1.6100 3.6600 1.8200 ;
        RECT 4.0600 1.6100 4.1800 1.8200 ;
        RECT 0.4200 0.4850 0.5400 0.7100 ;
        RECT 0.9400 0.4850 1.0600 0.7100 ;
        RECT 1.4600 0.4850 1.5800 0.7100 ;
        RECT 1.9800 0.4850 2.1000 0.7100 ;
        RECT 2.5000 0.4850 2.6200 0.7100 ;
        RECT 3.0200 0.4850 3.1400 0.7100 ;
        RECT 3.5400 0.4850 3.6600 0.7100 ;
        RECT 4.0600 0.4850 4.1800 0.7100 ;
    END
    ANTENNADIFFAREA 2.6 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 2.9000 1.1500 ;
    END
    ANTENNAGATEAREA 1.56 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.1700 1.7700 0.2700 2.0800 ;
        RECT 0.6900 1.7700 0.7900 2.0800 ;
        RECT 1.2100 1.7700 1.3100 2.0800 ;
        RECT 1.7300 1.7700 1.8300 2.0800 ;
        RECT 2.2500 1.7700 2.3500 2.0800 ;
        RECT 2.7700 1.7700 2.8700 2.0800 ;
        RECT 3.2900 1.7700 3.3900 2.0800 ;
        RECT 3.8100 1.7700 3.9100 2.0800 ;
        RECT 4.3300 1.7700 4.4300 2.0800 ;
    END
  END VDD
END INV_X16M_A12TH

MACRO INV_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.1450 0.3200 0.2450 0.8650 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 0.9850 0.1600 1.4050 ;
    END
    ANTENNAGATEAREA 0.0819 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 1.2900 0.5500 1.3900 ;
        RECT 0.4150 1.3900 0.5150 1.7200 ;
        RECT 0.4500 0.9100 0.5500 1.2900 ;
        RECT 0.4050 0.8100 0.5500 0.9100 ;
        RECT 0.4050 0.4600 0.5050 0.8100 ;
    END
    ANTENNADIFFAREA 0.238875 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.1450 1.7700 0.2450 2.0800 ;
    END
  END VDD
END INV_X1B_A12TH

MACRO INV_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9850 0.1600 1.4050 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9450 0.5500 1.2900 ;
        RECT 0.3500 1.2900 0.5500 1.3900 ;
        RECT 0.3500 0.8450 0.5500 0.9450 ;
        RECT 0.3500 1.3900 0.4500 1.7200 ;
        RECT 0.3500 0.4900 0.4500 0.8450 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.0850 1.7700 0.1950 2.0800 ;
    END
  END VDD
END INV_X1M_A12TH

MACRO INV_X1P2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7000 ;
        RECT 0.6150 0.3200 0.7150 0.7000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9500 0.7500 1.2500 ;
        RECT 0.3500 1.2500 0.7500 1.3500 ;
        RECT 0.3500 0.8500 0.7500 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7900 ;
        RECT 0.3500 0.5500 0.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0500 0.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.0972 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.4900 0.1900 2.0800 ;
        RECT 0.6100 1.4900 0.7100 2.0800 ;
    END
  END VDD
END INV_X1P2B_A12TH

MACRO INV_X1P2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.7750 ;
        RECT 0.6050 0.3200 0.7050 0.7050 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.0450 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1158 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.4500 0.7500 1.5500 ;
        RECT 0.3450 1.5500 0.4450 1.9600 ;
        RECT 0.6500 0.9000 0.7500 1.4500 ;
        RECT 0.3450 0.8000 0.7500 0.9000 ;
        RECT 0.3450 0.4200 0.4450 0.8000 ;
    END
    ANTENNADIFFAREA 0.193 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6050 1.6800 0.7050 2.0800 ;
        RECT 0.0850 1.6450 0.1850 2.0800 ;
    END
  END VDD
END INV_X1P2M_A12TH

MACRO INV_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7000 ;
        RECT 0.6100 0.3200 0.7100 0.7000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9500 0.7500 1.2500 ;
        RECT 0.3500 1.2500 0.7500 1.3500 ;
        RECT 0.3500 0.8500 0.7500 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7200 ;
        RECT 0.3500 0.6050 0.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0500 0.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.5050 0.1900 2.0800 ;
        RECT 0.6100 1.5050 0.7100 2.0800 ;
    END
  END VDD
END INV_X1P4B_A12TH

MACRO INV_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.8300 ;
        RECT 0.6050 0.3200 0.7050 0.7600 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 1.0500 0.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.4500 0.7500 1.5500 ;
        RECT 0.3450 1.5500 0.4450 1.8800 ;
        RECT 0.6500 0.9500 0.7500 1.4500 ;
        RECT 0.3450 0.8500 0.7500 0.9500 ;
        RECT 0.3450 0.4800 0.4450 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6050 1.6400 0.7050 2.0800 ;
        RECT 0.0850 1.6250 0.1850 2.0800 ;
    END
  END VDD
END INV_X1P4M_A12TH

MACRO INV_X1P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.8300 ;
        RECT 0.5750 0.3200 0.7450 0.7250 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9450 0.7500 1.2500 ;
        RECT 0.3500 1.2500 0.7500 1.3500 ;
        RECT 0.3500 0.8450 0.7500 0.9450 ;
        RECT 0.3500 1.3500 0.4500 1.7350 ;
        RECT 0.3500 0.4400 0.4500 0.8450 ;
    END
    ANTENNADIFFAREA 0.23 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.6800 0.1900 2.0800 ;
        RECT 0.6100 1.6300 0.7100 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1100 1.0500 0.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.138 ;
  END A
END INV_X1P7B_A12TH

MACRO INV_X1P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.7500 ;
        RECT 0.6050 0.3200 0.7050 0.7400 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 1.0500 0.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1638 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.4500 0.7500 1.5500 ;
        RECT 0.3450 1.5500 0.4450 1.8800 ;
        RECT 0.6500 0.9500 0.7500 1.4500 ;
        RECT 0.3450 0.8500 0.7500 0.9500 ;
        RECT 0.3450 0.4900 0.4450 0.8500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.6050 1.6600 0.7050 2.0800 ;
        RECT 0.0850 1.6250 0.1850 2.0800 ;
    END
  END VDD
END INV_X1P7M_A12TH

MACRO INV_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.8250 ;
        RECT 0.5750 0.3200 0.7450 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9500 0.7500 1.2500 ;
        RECT 0.3500 1.2500 0.7500 1.3500 ;
        RECT 0.3500 0.8500 0.7500 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7300 ;
        RECT 0.3500 0.4400 0.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6150 1.7700 0.7150 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1100 1.0500 0.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1638 ;
  END A
END INV_X2B_A12TH

MACRO INV_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.6500 ;
        RECT 0.6050 0.3200 0.7050 0.6500 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0500 0.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.195 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.4500 0.7500 1.5500 ;
        RECT 0.3450 1.5500 0.4450 1.8800 ;
        RECT 0.6500 0.9200 0.7500 1.4500 ;
        RECT 0.3450 0.8200 0.7500 0.9200 ;
        RECT 0.3450 0.5100 0.4450 0.8200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0850 1.7700 0.1850 2.0800 ;
        RECT 0.6050 1.7700 0.7050 2.0800 ;
    END
  END VDD
END INV_X2M_A12TH

MACRO INV_X2P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.1550 0.3200 0.2550 0.8450 ;
        RECT 0.6400 0.3200 0.8100 0.7400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.4150 1.2500 1.1500 1.3500 ;
        RECT 0.4150 0.8500 1.1500 0.9500 ;
        RECT 0.4150 1.3500 0.5150 1.7200 ;
        RECT 0.9350 1.3500 1.0350 1.7200 ;
        RECT 0.4150 0.4400 0.5150 0.8500 ;
        RECT 0.9350 0.4400 1.0350 0.8500 ;
    END
    ANTENNADIFFAREA 0.4617 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.6750 1.6300 0.7750 2.0800 ;
        RECT 0.1550 1.6200 0.2550 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3100 1.0500 0.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.2052 ;
  END A
END INV_X2P5B_A12TH

MACRO INV_X2P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.1600 0.3200 0.2600 0.7100 ;
        RECT 0.6800 0.3200 0.7800 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.4200 1.2500 1.1500 1.3500 ;
        RECT 0.4200 0.8500 1.1500 0.9500 ;
        RECT 0.4200 1.3500 0.5200 1.7200 ;
        RECT 0.9400 1.3500 1.0400 1.7200 ;
        RECT 0.4200 0.4500 0.5200 0.8500 ;
        RECT 0.9400 0.4500 1.0400 0.8500 ;
    END
    ANTENNADIFFAREA 0.51 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 0.8250 1.1500 ;
    END
    ANTENNAGATEAREA 0.2448 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.1550 1.6200 0.2650 2.0800 ;
        RECT 0.6750 1.6200 0.7850 2.0800 ;
    END
  END VDD
END INV_X2P5M_A12TH

MACRO FILLTIE16_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.5150 1.9900 0.6850 2.0800 ;
        RECT 0.9200 1.9900 1.0900 2.0800 ;
        RECT 1.3200 1.9900 1.4900 2.0800 ;
        RECT 1.7200 1.9900 1.8900 2.0800 ;
        RECT 2.1200 1.9900 2.2900 2.0800 ;
        RECT 2.5200 1.9900 2.6900 2.0800 ;
        RECT 0.1500 1.5050 0.2500 2.0800 ;
        RECT 2.9500 1.5050 3.0500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1500 0.3200 0.2500 0.8550 ;
        RECT 0.5150 0.3200 0.6850 0.4100 ;
        RECT 0.9150 0.3200 1.0850 0.4100 ;
        RECT 1.3150 0.3200 1.4850 0.4100 ;
        RECT 1.7150 0.3200 1.8850 0.4100 ;
        RECT 2.1150 0.3200 2.2850 0.4100 ;
        RECT 2.5150 0.3200 2.6850 0.4100 ;
        RECT 2.9500 0.3200 3.0500 0.8550 ;
    END
  END VSS
END FILLTIE16_A12TH

MACRO FILLTIE2_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.4450 2.7200 ;
        RECT 0.1500 1.4500 0.2500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.4450 0.3200 ;
        RECT 0.1500 0.3200 0.2500 0.8450 ;
    END
  END VSS
END FILLTIE2_A12TH

MACRO FILLTIE32_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.5150 1.9900 0.6850 2.0800 ;
        RECT 0.9200 1.9900 1.0900 2.0800 ;
        RECT 1.3200 1.9900 1.4900 2.0800 ;
        RECT 1.7200 1.9900 1.8900 2.0800 ;
        RECT 2.1200 1.9900 2.2900 2.0800 ;
        RECT 2.5200 1.9900 2.6900 2.0800 ;
        RECT 2.9150 1.9900 3.0850 2.0800 ;
        RECT 3.3200 1.9900 3.4900 2.0800 ;
        RECT 3.7200 1.9900 3.8900 2.0800 ;
        RECT 4.1200 1.9900 4.2900 2.0800 ;
        RECT 4.5200 1.9900 4.6900 2.0800 ;
        RECT 4.9200 1.9900 5.0900 2.0800 ;
        RECT 5.3200 1.9900 5.4900 2.0800 ;
        RECT 5.7200 1.9900 5.8900 2.0800 ;
        RECT 0.1500 1.5050 0.2500 2.0800 ;
        RECT 6.1500 1.5050 6.2500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.1500 0.3200 0.2500 0.8550 ;
        RECT 0.5150 0.3200 0.6850 0.4100 ;
        RECT 0.9150 0.3200 1.0850 0.4100 ;
        RECT 1.3150 0.3200 1.4850 0.4100 ;
        RECT 1.7150 0.3200 1.8850 0.4100 ;
        RECT 2.1150 0.3200 2.2850 0.4100 ;
        RECT 2.5150 0.3200 2.6850 0.4100 ;
        RECT 2.9150 0.3200 3.0850 0.4100 ;
        RECT 3.3150 0.3200 3.4850 0.4100 ;
        RECT 3.7150 0.3200 3.8850 0.4100 ;
        RECT 4.1150 0.3200 4.2850 0.4100 ;
        RECT 4.5150 0.3200 4.6850 0.4100 ;
        RECT 4.9150 0.3200 5.0850 0.4100 ;
        RECT 5.3150 0.3200 5.4850 0.4100 ;
        RECT 5.7150 0.3200 5.8850 0.4100 ;
        RECT 6.1500 0.3200 6.2500 0.8550 ;
    END
  END VSS
END FILLTIE32_A12TH

MACRO FILLTIE4_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.1350 1.4500 0.2350 2.0800 ;
        RECT 0.5250 1.4500 0.6250 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.8550 ;
        RECT 0.5150 0.3200 0.6150 0.8550 ;
    END
  END VSS
END FILLTIE4_A12TH

MACRO FILLTIE64_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.8450 2.7200 ;
        RECT 0.5150 1.9900 0.6850 2.0800 ;
        RECT 0.9200 1.9900 1.0900 2.0800 ;
        RECT 1.3200 1.9900 1.4900 2.0800 ;
        RECT 1.7200 1.9900 1.8900 2.0800 ;
        RECT 2.1200 1.9900 2.2900 2.0800 ;
        RECT 2.5200 1.9900 2.6900 2.0800 ;
        RECT 2.9150 1.9900 3.0850 2.0800 ;
        RECT 3.3200 1.9900 3.4900 2.0800 ;
        RECT 3.7200 1.9900 3.8900 2.0800 ;
        RECT 4.1200 1.9900 4.2900 2.0800 ;
        RECT 4.5200 1.9900 4.6900 2.0800 ;
        RECT 4.9200 1.9900 5.0900 2.0800 ;
        RECT 5.3200 1.9900 5.4900 2.0800 ;
        RECT 5.7200 1.9900 5.8900 2.0800 ;
        RECT 6.1150 1.9900 6.2850 2.0800 ;
        RECT 6.5200 1.9900 6.6900 2.0800 ;
        RECT 6.9200 1.9900 7.0900 2.0800 ;
        RECT 7.3200 1.9900 7.4900 2.0800 ;
        RECT 7.7200 1.9900 7.8900 2.0800 ;
        RECT 8.1200 1.9900 8.2900 2.0800 ;
        RECT 8.5150 1.9900 8.6850 2.0800 ;
        RECT 8.9200 1.9900 9.0900 2.0800 ;
        RECT 9.3200 1.9900 9.4900 2.0800 ;
        RECT 9.7200 1.9900 9.8900 2.0800 ;
        RECT 10.1200 1.9900 10.2900 2.0800 ;
        RECT 10.5200 1.9900 10.6900 2.0800 ;
        RECT 10.9200 1.9900 11.0900 2.0800 ;
        RECT 11.3200 1.9900 11.4900 2.0800 ;
        RECT 11.7200 1.9900 11.8900 2.0800 ;
        RECT 12.1200 1.9900 12.2900 2.0800 ;
        RECT 0.1500 1.5050 0.2500 2.0800 ;
        RECT 12.5500 1.5050 12.6500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.8450 0.3200 ;
        RECT 0.1500 0.3200 0.2500 0.8550 ;
        RECT 0.5150 0.3200 0.6850 0.4100 ;
        RECT 0.9150 0.3200 1.0850 0.4100 ;
        RECT 1.3150 0.3200 1.4850 0.4100 ;
        RECT 1.7150 0.3200 1.8850 0.4100 ;
        RECT 2.1150 0.3200 2.2850 0.4100 ;
        RECT 2.5150 0.3200 2.6850 0.4100 ;
        RECT 2.9150 0.3200 3.0850 0.4100 ;
        RECT 3.3150 0.3200 3.4850 0.4100 ;
        RECT 3.7150 0.3200 3.8850 0.4100 ;
        RECT 4.1150 0.3200 4.2850 0.4100 ;
        RECT 4.5150 0.3200 4.6850 0.4100 ;
        RECT 4.9150 0.3200 5.0850 0.4100 ;
        RECT 5.3150 0.3200 5.4850 0.4100 ;
        RECT 5.7150 0.3200 5.8850 0.4100 ;
        RECT 6.1150 0.3200 6.2850 0.4100 ;
        RECT 6.5150 0.3200 6.6850 0.4100 ;
        RECT 6.9150 0.3200 7.0850 0.4100 ;
        RECT 7.3150 0.3200 7.4850 0.4100 ;
        RECT 7.7150 0.3200 7.8850 0.4100 ;
        RECT 8.1150 0.3200 8.2850 0.4100 ;
        RECT 8.5150 0.3200 8.6850 0.4100 ;
        RECT 8.9150 0.3200 9.0850 0.4100 ;
        RECT 9.3150 0.3200 9.4850 0.4100 ;
        RECT 9.7150 0.3200 9.8850 0.4100 ;
        RECT 10.1150 0.3200 10.2850 0.4100 ;
        RECT 10.5150 0.3200 10.6850 0.4100 ;
        RECT 10.9150 0.3200 11.0850 0.4100 ;
        RECT 11.3150 0.3200 11.4850 0.4100 ;
        RECT 11.7150 0.3200 11.8850 0.4100 ;
        RECT 12.1150 0.3200 12.2850 0.4100 ;
        RECT 12.5550 0.3200 12.6550 0.8550 ;
    END
  END VSS
END FILLTIE64_A12TH

MACRO FILLTIE8_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.5150 1.9900 0.6850 2.0800 ;
        RECT 0.9150 1.9900 1.0850 2.0800 ;
        RECT 0.1350 1.5050 0.2350 2.0800 ;
        RECT 1.3500 1.5050 1.4500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.8550 ;
        RECT 0.5150 0.3200 0.6850 0.4100 ;
        RECT 0.9150 0.3200 1.0850 0.4100 ;
        RECT 1.3500 0.3200 1.4500 0.8550 ;
    END
  END VSS
END FILLTIE8_A12TH

MACRO FRICG_X0P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9050 ;
        RECT 1.1350 0.3200 1.2250 0.8750 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8300 1.5500 1.5250 ;
        RECT 1.3950 1.5250 1.5500 1.6250 ;
        RECT 1.3350 0.7300 1.5500 0.8300 ;
        RECT 1.3950 1.6250 1.4950 1.9550 ;
    END
    ANTENNADIFFAREA 0.111075 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1300 1.5550 1.2200 2.0800 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6800 0.1700 1.4100 ;
      RECT 0.3400 1.3000 0.7500 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7150 ;
      RECT 0.8600 1.3050 1.3300 1.3950 ;
      RECT 1.2400 1.0750 1.3300 1.3050 ;
      RECT 0.9500 0.9850 1.3300 1.0750 ;
      RECT 0.8600 1.3950 0.9500 1.7150 ;
      RECT 0.9500 0.8250 1.0400 0.9850 ;
      RECT 0.8000 0.7350 1.0400 0.8250 ;
  END
END FRICG_X0P5B_A12TH

MACRO FRICG_X0P6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9050 ;
        RECT 1.1350 0.3200 1.2250 0.8500 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8550 1.5500 1.5250 ;
        RECT 1.3950 1.5250 1.5500 1.6250 ;
        RECT 1.3350 0.7550 1.5500 0.8550 ;
        RECT 1.3950 1.6250 1.4950 1.9550 ;
    END
    ANTENNADIFFAREA 0.133125 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1200 1.5550 1.2100 2.0800 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6800 0.1700 1.4100 ;
      RECT 0.3400 1.2950 0.7250 1.3850 ;
      RECT 0.3400 1.3850 0.4300 1.7150 ;
      RECT 0.8600 1.3100 1.3300 1.4000 ;
      RECT 1.2400 1.0600 1.3300 1.3100 ;
      RECT 0.9500 0.9700 1.3300 1.0600 ;
      RECT 0.8600 1.4000 0.9500 1.7150 ;
      RECT 0.9500 0.8250 1.0400 0.9700 ;
      RECT 0.8000 0.7350 1.0400 0.8250 ;
  END
END FRICG_X0P6B_A12TH

MACRO FRICG_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9050 ;
        RECT 1.1350 0.3200 1.2250 0.8500 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9050 1.5500 1.5250 ;
        RECT 1.3950 1.5250 1.5500 1.6250 ;
        RECT 1.3350 0.8050 1.5500 0.9050 ;
        RECT 1.3950 1.6250 1.4950 1.9550 ;
    END
    ANTENNADIFFAREA 0.155975 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1350 1.5550 1.2250 2.0800 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6800 0.1700 1.4100 ;
      RECT 0.3400 1.3000 0.8250 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7150 ;
      RECT 0.9500 1.2850 1.3300 1.3750 ;
      RECT 1.2400 1.1250 1.3300 1.2850 ;
      RECT 0.8000 1.5650 1.0400 1.6550 ;
      RECT 0.9500 1.3750 1.0400 1.5650 ;
      RECT 0.9500 0.8150 1.0400 1.2850 ;
      RECT 0.8000 0.7250 1.0400 0.8150 ;
  END
END FRICG_X0P7B_A12TH

MACRO FRICG_X0P8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9050 ;
        RECT 1.1350 0.3200 1.2250 0.9850 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9950 1.5500 1.4100 ;
        RECT 1.3950 1.4100 1.5500 1.5100 ;
        RECT 1.3900 0.8950 1.5500 0.9950 ;
        RECT 1.3950 1.5100 1.4950 1.8400 ;
        RECT 1.3900 0.5850 1.4900 0.8950 ;
    END
    ANTENNADIFFAREA 0.17805 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1350 1.6050 1.2250 2.0800 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6800 0.1700 1.4100 ;
      RECT 0.3400 1.3000 0.8250 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7150 ;
      RECT 0.9500 1.1500 1.3400 1.2500 ;
      RECT 0.8000 1.5650 1.0400 1.6550 ;
      RECT 0.9500 1.2500 1.0400 1.5650 ;
      RECT 0.9500 0.8150 1.0400 1.1500 ;
      RECT 0.8000 0.7250 1.0400 0.8150 ;
  END
END FRICG_X0P8B_A12TH

MACRO FRICG_X11B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9700 ;
        RECT 1.3750 0.3200 1.4650 0.6600 ;
        RECT 2.3700 0.3200 2.4600 0.6600 ;
        RECT 2.9200 0.3200 3.0100 0.5100 ;
        RECT 3.4400 0.3200 3.5300 0.5100 ;
        RECT 3.9600 0.3200 4.0500 0.5100 ;
        RECT 4.4800 0.3200 4.5700 0.5100 ;
        RECT 5.0000 0.3200 5.0900 0.7300 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6200 0.8600 4.7800 1.2200 ;
        RECT 2.6550 1.2200 4.8400 1.3800 ;
        RECT 2.6550 0.7000 4.8350 0.8600 ;
        RECT 2.6550 1.3800 2.7550 1.7250 ;
        RECT 3.1750 1.3800 3.2750 1.7250 ;
        RECT 3.6950 1.3800 3.7950 1.7250 ;
        RECT 4.2150 1.3800 4.3150 1.7250 ;
        RECT 4.7300 1.3800 4.8400 1.7250 ;
        RECT 2.6550 0.4150 2.7550 0.7000 ;
        RECT 3.1750 0.4150 3.2750 0.7000 ;
        RECT 3.6950 0.4150 3.7950 0.7000 ;
        RECT 4.2150 0.4150 4.3150 0.7000 ;
        RECT 4.7350 0.4150 4.8350 0.7000 ;
    END
    ANTENNADIFFAREA 1.6146 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0550 1.2750 2.0900 1.3500 ;
        RECT 0.7500 1.2500 2.0900 1.2750 ;
        RECT 0.7500 1.1750 1.1550 1.2500 ;
    END
    ANTENNAGATEAREA 0.3432 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 0.6750 1.8850 0.7650 2.0800 ;
        RECT 2.9200 1.7700 3.0100 2.0800 ;
        RECT 3.4400 1.7700 3.5300 2.0800 ;
        RECT 3.9600 1.7700 4.0500 2.0800 ;
        RECT 4.4800 1.7700 4.5700 2.0800 ;
        RECT 5.0000 1.7700 5.0900 2.0800 ;
        RECT 1.7500 1.7650 1.8400 2.0800 ;
        RECT 1.1950 1.6850 1.2850 2.0800 ;
        RECT 0.0800 1.6450 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.2450 0.2300 1.4150 ;
      RECT 0.0800 0.7650 0.1700 1.2450 ;
      RECT 0.5500 0.9950 2.3100 1.0850 ;
      RECT 1.2600 1.0850 1.5800 1.1450 ;
      RECT 2.2200 1.0850 2.3100 1.2550 ;
      RECT 0.3400 1.3750 0.4300 1.6700 ;
      RECT 0.3400 1.2850 0.6400 1.3750 ;
      RECT 0.5500 1.0850 0.6400 1.2850 ;
      RECT 2.4350 0.9750 4.3650 1.0650 ;
      RECT 0.9350 1.5750 1.0250 1.9350 ;
      RECT 0.9150 0.4450 1.0050 0.7850 ;
      RECT 1.4450 1.5750 1.5350 1.9350 ;
      RECT 2.0100 1.5750 2.1000 1.9350 ;
      RECT 1.8350 0.4450 1.9250 0.7850 ;
      RECT 0.9350 1.4850 2.5250 1.5750 ;
      RECT 2.4350 1.0650 2.5250 1.4850 ;
      RECT 2.4350 0.8750 2.5250 0.9750 ;
      RECT 0.9150 0.7850 2.5250 0.8750 ;
  END
END FRICG_X11B_A12TH

MACRO FRICG_X13B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9050 ;
        RECT 1.3750 0.3200 1.4650 0.6300 ;
        RECT 2.3250 0.3200 2.4150 0.6300 ;
        RECT 3.0750 0.3200 3.1650 0.7500 ;
        RECT 3.5550 0.3200 3.7250 0.6900 ;
        RECT 4.0750 0.3200 4.2450 0.6900 ;
        RECT 4.5950 0.3200 4.7650 0.6900 ;
        RECT 5.1150 0.3200 5.2850 0.6900 ;
        RECT 5.6350 0.3200 5.8050 0.6900 ;
        RECT 6.1550 0.3200 6.3250 0.6900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.1500 1.1500 ;
        RECT 1.0500 1.0350 1.1500 1.0500 ;
        RECT 1.0500 0.9350 1.8300 1.0350 ;
        RECT 1.7300 1.0350 1.8300 1.0500 ;
        RECT 1.7300 1.0500 2.8000 1.1500 ;
        RECT 2.7000 1.1500 2.8000 1.2650 ;
    END
    ANTENNAGATEAREA 0.405 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8100 0.9600 6.0300 1.4100 ;
        RECT 3.0750 1.4100 6.2900 1.5900 ;
        RECT 3.3300 0.7800 6.0300 0.9600 ;
        RECT 3.0750 1.5900 3.1650 1.8500 ;
        RECT 3.5900 1.5900 3.6900 1.8500 ;
        RECT 4.1100 1.5900 4.2100 1.8500 ;
        RECT 4.6300 1.5900 4.7300 1.8500 ;
        RECT 5.1500 1.5900 5.2500 1.8500 ;
        RECT 5.6700 1.5900 5.7700 1.8500 ;
        RECT 6.1900 1.5900 6.2900 1.8500 ;
        RECT 3.3300 0.4100 3.4300 0.7800 ;
        RECT 3.8500 0.4100 3.9500 0.7800 ;
        RECT 4.3700 0.4100 4.4700 0.7800 ;
        RECT 4.8900 0.4100 4.9900 0.7800 ;
        RECT 5.4100 0.4100 5.5100 0.7800 ;
        RECT 5.9300 0.4100 6.0300 0.7800 ;
    END
    ANTENNADIFFAREA 1.9396 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.6750 1.9100 0.7650 2.0800 ;
        RECT 1.5300 1.7700 1.6200 2.0800 ;
        RECT 2.0950 1.7700 2.1850 2.0800 ;
        RECT 2.8150 1.7700 2.9050 2.0800 ;
        RECT 3.3350 1.7700 3.4250 2.0800 ;
        RECT 3.8550 1.7700 3.9450 2.0800 ;
        RECT 4.3750 1.7700 4.4650 2.0800 ;
        RECT 4.8950 1.7700 4.9850 2.0800 ;
        RECT 5.4150 1.7700 5.5050 2.0800 ;
        RECT 5.9350 1.7700 6.0250 2.0800 ;
        RECT 1.1950 1.7400 1.2850 2.0800 ;
        RECT 0.0800 1.6950 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6950 0.1700 1.3600 ;
      RECT 0.3400 1.4200 0.4300 1.6300 ;
      RECT 0.3400 1.3300 2.5500 1.4200 ;
      RECT 0.4700 1.0500 0.5600 1.3300 ;
      RECT 1.2400 1.1650 1.6100 1.4200 ;
      RECT 2.8950 1.0700 5.4800 1.1600 ;
      RECT 0.9350 1.6400 1.0250 1.9800 ;
      RECT 0.9150 0.4300 1.0050 0.7500 ;
      RECT 1.8350 1.6400 1.9250 1.9800 ;
      RECT 1.8350 0.4300 1.9250 0.7500 ;
      RECT 2.5400 1.6400 2.6300 1.9800 ;
      RECT 0.9350 1.5500 2.9850 1.6400 ;
      RECT 2.8950 1.1600 2.9850 1.5500 ;
      RECT 2.8950 0.8400 2.9850 1.0700 ;
      RECT 0.9150 0.7500 2.9850 0.8400 ;
      RECT 2.8250 0.4250 2.9150 0.7500 ;
  END
END FRICG_X13B_A12TH

MACRO FRICG_X16B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.6500 ;
        RECT 1.3750 0.3200 1.4650 0.6300 ;
        RECT 2.3250 0.3200 2.4150 0.6300 ;
        RECT 3.1900 0.3200 3.2800 0.8000 ;
        RECT 3.7100 0.3200 3.8000 0.5800 ;
        RECT 4.2300 0.3200 4.3200 0.5800 ;
        RECT 4.7500 0.3200 4.8400 0.5800 ;
        RECT 5.2700 0.3200 5.3600 0.5800 ;
        RECT 5.7900 0.3200 5.8800 0.5800 ;
        RECT 6.3100 0.3200 6.4000 0.5800 ;
        RECT 6.8300 0.3200 6.9200 0.5800 ;
        RECT 7.3500 0.3200 7.4400 0.8000 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9900 0.9250 7.2100 1.2900 ;
        RECT 3.4500 1.2900 7.2100 1.5100 ;
        RECT 3.4500 0.7050 7.2100 0.9250 ;
        RECT 3.4500 1.5100 3.5400 1.7200 ;
        RECT 3.9700 1.5100 4.0600 1.7200 ;
        RECT 4.4900 1.5100 4.5800 1.7200 ;
        RECT 5.0100 1.5100 5.1000 1.7200 ;
        RECT 5.5300 1.5100 5.6200 1.7200 ;
        RECT 6.0500 1.5100 6.1400 1.7200 ;
        RECT 6.5700 1.5100 6.6600 1.7200 ;
        RECT 7.0800 1.5100 7.2100 1.7200 ;
        RECT 3.4500 0.4150 3.5400 0.7050 ;
        RECT 3.9700 0.4150 4.0600 0.7050 ;
        RECT 4.4900 0.4150 4.5800 0.7050 ;
        RECT 5.0100 0.4150 5.1000 0.7050 ;
        RECT 5.5300 0.4150 5.6200 0.7050 ;
        RECT 6.0500 0.4150 6.1400 0.7050 ;
        RECT 6.5700 0.4150 6.6600 0.7050 ;
        RECT 7.0800 0.4150 7.2100 0.7050 ;
    END
    ANTENNADIFFAREA 2.376 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7450 1.0500 1.1500 1.2200 ;
        RECT 1.0500 1.0450 1.1500 1.0500 ;
        RECT 1.0500 0.9450 1.8150 1.0450 ;
        RECT 1.7150 1.0450 1.8150 1.0500 ;
        RECT 1.7150 1.0500 2.1050 1.2400 ;
        RECT 2.0050 1.0350 2.1050 1.0500 ;
        RECT 2.0050 0.9350 2.8100 1.0350 ;
        RECT 2.7100 1.0350 2.8100 1.3100 ;
    END
    ANTENNAGATEAREA 0.495 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.6450 2.7200 ;
        RECT 0.6750 1.7700 0.7650 2.0800 ;
        RECT 1.1950 1.7700 1.2850 2.0800 ;
        RECT 1.5300 1.7700 1.6200 2.0800 ;
        RECT 2.0950 1.7700 2.1850 2.0800 ;
        RECT 2.8150 1.7700 2.9050 2.0800 ;
        RECT 3.1900 1.7700 3.2800 2.0800 ;
        RECT 3.7100 1.7700 3.8000 2.0800 ;
        RECT 4.2300 1.7700 4.3200 2.0800 ;
        RECT 4.7500 1.7700 4.8400 2.0800 ;
        RECT 5.2700 1.7700 5.3600 2.0800 ;
        RECT 5.7900 1.7700 5.8800 2.0800 ;
        RECT 6.3100 1.7700 6.4000 2.0800 ;
        RECT 6.8300 1.7700 6.9200 2.0800 ;
        RECT 7.3500 1.7700 7.4400 2.0800 ;
        RECT 0.0800 1.7650 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.9500 1.0700 6.5250 1.1600 ;
      RECT 0.9350 1.5500 3.0400 1.6400 ;
      RECT 2.9500 1.1600 3.0400 1.5500 ;
      RECT 2.9500 0.8400 3.0400 1.0700 ;
      RECT 0.8600 0.7500 3.0400 0.8400 ;
      RECT 2.8250 0.4100 2.9150 0.7500 ;
      RECT 0.9350 1.6400 1.0250 1.9800 ;
      RECT 0.8600 0.4100 0.9500 0.7500 ;
      RECT 1.8350 1.6400 1.9250 1.9800 ;
      RECT 1.8350 0.4100 1.9250 0.7500 ;
      RECT 2.5400 1.6400 2.6300 1.9800 ;
      RECT 0.0800 0.4400 0.1700 1.2950 ;
      RECT 0.3400 1.4250 0.4300 1.5550 ;
      RECT 0.3400 1.3350 2.3000 1.4250 ;
      RECT 0.4750 1.0850 0.5650 1.3350 ;
      RECT 2.2100 1.2350 2.3000 1.3350 ;
      RECT 2.2100 1.1450 2.5800 1.2350 ;
      RECT 1.2400 1.1650 1.6100 1.4250 ;
  END
END FRICG_X16B_A12TH

MACRO FRICG_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.8900 ;
        RECT 1.1350 0.3200 1.2250 0.8950 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
        RECT 1.1350 1.4950 1.2250 2.0800 ;
    END
  END VDD

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9200 1.5500 1.3250 ;
        RECT 1.3950 1.3250 1.5500 1.4250 ;
        RECT 1.3900 0.8200 1.5500 0.9200 ;
        RECT 1.3950 1.4250 1.4950 1.7550 ;
        RECT 1.3900 0.4900 1.4900 0.8200 ;
    END
    ANTENNADIFFAREA 0.22295 ;
  END ECK
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6650 0.1700 1.4100 ;
      RECT 0.3400 1.3000 0.8250 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7150 ;
      RECT 0.9500 1.1300 1.3300 1.2200 ;
      RECT 1.2400 1.0100 1.3300 1.1300 ;
      RECT 0.8000 1.5650 1.0400 1.6550 ;
      RECT 0.9500 1.2200 1.0400 1.5650 ;
      RECT 0.9500 0.6850 1.0400 1.1300 ;
      RECT 0.8300 0.5950 1.0400 0.6850 ;
  END
END FRICG_X1B_A12TH

MACRO FRICG_X1P2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.8700 ;
        RECT 1.1950 0.3200 1.2850 0.9050 ;
        RECT 1.7150 0.3200 1.8050 0.9050 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7600 1.5500 1.8200 ;
    END
    ANTENNADIFFAREA 0.165 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.1950 1.5100 1.2850 2.0800 ;
        RECT 1.7150 1.5100 1.8050 2.0800 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6600 0.1700 1.4100 ;
      RECT 0.3400 1.3000 0.8250 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7150 ;
      RECT 0.9500 1.2150 1.3400 1.3050 ;
      RECT 1.2500 1.0950 1.3400 1.2150 ;
      RECT 0.8000 1.5650 1.0400 1.6550 ;
      RECT 0.9500 1.3050 1.0400 1.5650 ;
      RECT 0.9500 0.8650 1.0400 1.2150 ;
      RECT 0.8950 0.7750 1.0400 0.8650 ;
      RECT 0.8950 0.4600 0.9850 0.7750 ;
  END
END FRICG_X1P2B_A12TH

MACRO FRICG_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3750 0.3200 0.4650 0.8800 ;
        RECT 1.1950 0.3200 1.2850 0.8800 ;
        RECT 1.7150 0.3200 1.8050 0.9850 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7600 1.5500 1.7950 ;
    END
    ANTENNADIFFAREA 0.194025 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4350 1.0500 0.8550 1.1500 ;
    END
    ANTENNAGATEAREA 0.0516 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.1950 1.5850 1.2850 2.0800 ;
        RECT 1.7150 1.5850 1.8050 2.0800 ;
        RECT 0.0800 1.5050 0.1700 2.0800 ;
        RECT 0.6000 1.5050 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6550 0.1700 1.4100 ;
      RECT 0.3400 1.3000 0.8250 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7150 ;
      RECT 0.9550 1.1250 1.3500 1.2150 ;
      RECT 0.8000 1.5650 1.0450 1.6550 ;
      RECT 0.9550 1.2150 1.0450 1.5650 ;
      RECT 0.9550 0.8750 1.0450 1.1250 ;
      RECT 0.8950 0.7850 1.0450 0.8750 ;
      RECT 0.8950 0.4400 0.9850 0.7850 ;
  END
END FRICG_X1P4B_A12TH

MACRO FRICG_X1P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3750 0.3200 0.4650 0.8700 ;
        RECT 1.1950 0.3200 1.2850 0.9450 ;
        RECT 1.7150 0.3200 1.8050 0.9750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4200 1.0500 0.8500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0606 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.5800 1.5500 1.7150 ;
    END
    ANTENNADIFFAREA 0.232 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.7150 1.6800 1.8050 2.0800 ;
        RECT 0.6000 1.6350 0.6900 2.0800 ;
        RECT 0.0800 1.6100 0.1700 2.0800 ;
        RECT 1.1950 1.3950 1.2850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6450 0.1700 1.4100 ;
      RECT 0.3400 1.4550 0.8200 1.5450 ;
      RECT 0.3400 1.5450 0.4300 1.8400 ;
      RECT 1.0050 1.1550 1.3600 1.2450 ;
      RECT 1.2700 1.0550 1.3600 1.1550 ;
      RECT 0.8000 1.6900 1.0950 1.7800 ;
      RECT 1.0050 1.2450 1.0950 1.6900 ;
      RECT 1.0050 0.8650 1.0950 1.1550 ;
      RECT 0.9150 0.7750 1.0950 0.8650 ;
      RECT 0.9150 0.4100 1.0050 0.7750 ;
  END
END FRICG_X1P7B_A12TH

MACRO FRICG_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9050 ;
        RECT 1.1950 0.3200 1.2850 0.9250 ;
        RECT 1.7150 0.3200 1.8050 0.9250 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.5200 1.5500 1.7000 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0500 0.8650 1.1500 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.1950 1.7700 1.2850 2.0800 ;
        RECT 1.7150 1.7700 1.8050 2.0800 ;
        RECT 0.6150 1.6900 0.7050 2.0800 ;
        RECT 0.0800 1.6550 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6800 0.1700 1.4100 ;
      RECT 0.3400 1.4550 0.8400 1.5450 ;
      RECT 0.3400 1.5450 0.4300 1.9000 ;
      RECT 0.9650 1.1450 1.3400 1.2350 ;
      RECT 1.2500 1.0350 1.3400 1.1450 ;
      RECT 0.8150 1.7500 1.0550 1.8400 ;
      RECT 0.9650 1.2350 1.0550 1.7500 ;
      RECT 0.9650 0.9000 1.0550 1.1450 ;
      RECT 0.8950 0.8100 1.0550 0.9000 ;
      RECT 0.8950 0.4450 0.9850 0.8100 ;
  END
END FRICG_X2B_A12TH

MACRO FRICG_X2P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.8950 ;
        RECT 1.2100 0.3200 1.3000 0.9600 ;
        RECT 1.7250 0.3200 1.8250 0.7500 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.6150 1.6900 0.7050 2.0800 ;
        RECT 0.0800 1.6600 0.1700 2.0800 ;
        RECT 1.2100 1.6200 1.3000 2.0800 ;
        RECT 1.7300 1.6200 1.8200 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0500 0.8650 1.1500 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.2500 ;
        RECT 1.4650 1.2500 2.0850 1.3500 ;
        RECT 1.4650 0.8500 2.0850 0.9500 ;
        RECT 1.4650 1.3500 1.5650 1.7200 ;
        RECT 1.9850 1.3500 2.0850 1.7200 ;
        RECT 1.4650 0.5500 1.5650 0.8500 ;
        RECT 1.9850 0.5300 2.0850 0.8500 ;
    END
    ANTENNADIFFAREA 0.415 ;
  END ECK
  OBS
    LAYER M1 ;
      RECT 0.0800 0.6700 0.1700 1.4100 ;
      RECT 0.3400 1.4550 0.8400 1.5450 ;
      RECT 0.3400 1.5450 0.4300 1.9000 ;
      RECT 0.9650 1.0550 1.7400 1.1450 ;
      RECT 0.8150 1.7500 1.0550 1.8400 ;
      RECT 0.9650 1.1450 1.0550 1.7500 ;
      RECT 0.9650 0.8900 1.0550 1.0550 ;
      RECT 0.8950 0.8000 1.0550 0.8900 ;
      RECT 0.8950 0.4550 0.9850 0.8000 ;
  END
END FRICG_X2P5B_A12TH

MACRO FRICG_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3950 0.3200 0.5650 0.5800 ;
        RECT 1.2450 0.3200 1.3350 0.9150 ;
        RECT 1.7650 0.3200 1.8550 0.6950 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 1.0500 0.8100 1.1500 ;
        RECT 0.7100 1.1500 0.8100 1.1600 ;
        RECT 0.7100 1.1600 0.9550 1.2600 ;
    END
    ANTENNAGATEAREA 0.1002 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.2500 ;
        RECT 1.5000 1.2500 2.1200 1.3500 ;
        RECT 1.5000 0.8500 2.1200 0.9500 ;
        RECT 1.5000 1.3500 1.6000 1.7200 ;
        RECT 2.0200 1.3500 2.1200 1.7200 ;
        RECT 2.0200 0.5100 2.1200 0.8500 ;
        RECT 1.5000 0.5050 1.6000 0.8500 ;
    END
    ANTENNADIFFAREA 0.53195 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.2050 1.7950 1.2950 2.0800 ;
        RECT 1.7650 1.7700 1.8550 2.0800 ;
        RECT 0.6150 1.6350 0.7050 2.0800 ;
        RECT 0.0800 1.6050 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7750 0.1700 1.5050 ;
      RECT 0.3400 1.4550 0.8400 1.5450 ;
      RECT 0.3400 1.5450 0.4300 1.8250 ;
      RECT 1.0550 1.0550 1.7350 1.1450 ;
      RECT 0.8750 1.7250 0.9650 1.8500 ;
      RECT 0.8750 1.6350 1.1450 1.7250 ;
      RECT 1.0550 1.1450 1.1450 1.6350 ;
      RECT 1.0550 0.9600 1.1450 1.0550 ;
      RECT 0.8950 0.8700 1.1450 0.9600 ;
      RECT 0.8950 0.5500 0.9850 0.8700 ;
  END
END FRICG_X3B_A12TH

MACRO FRICG_X3P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9550 ;
        RECT 1.3900 0.3200 1.4800 0.6550 ;
        RECT 1.8050 0.3200 1.8950 0.6500 ;
        RECT 2.2850 0.3200 2.4550 0.5500 ;
    END
  END VSS

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7500 2.7500 1.2500 ;
        RECT 2.0600 1.2500 2.7500 1.3500 ;
        RECT 2.0650 0.6500 2.7500 0.7500 ;
        RECT 2.0600 1.3500 2.1600 1.6800 ;
        RECT 2.5850 1.3500 2.6750 1.7200 ;
        RECT 2.0650 0.5200 2.1550 0.6500 ;
        RECT 2.5450 0.4100 2.7150 0.6500 ;
    END
    ANTENNADIFFAREA 0.57765 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.2100 1.7900 1.3000 2.0800 ;
        RECT 1.8050 1.7700 1.8950 2.0800 ;
        RECT 2.3250 1.7700 2.4150 2.0800 ;
        RECT 0.6900 1.5700 0.7800 2.0800 ;
        RECT 0.0800 1.5600 0.1700 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7100 1.0500 1.1400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1152 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7450 0.1700 1.4400 ;
      RECT 0.3400 1.3000 1.4650 1.3900 ;
      RECT 0.3400 1.3900 0.4300 1.7050 ;
      RECT 1.6100 0.9000 2.4550 0.9500 ;
      RECT 0.8550 0.8600 2.4550 0.9000 ;
      RECT 0.9500 1.6400 1.0400 1.9600 ;
      RECT 0.8550 0.4700 0.9450 0.8100 ;
      RECT 0.9500 1.5500 1.7000 1.6400 ;
      RECT 1.6100 0.9500 1.7000 1.5500 ;
      RECT 0.8550 0.8100 1.7000 0.8600 ;
  END
END FRICG_X3P5B_A12TH

MACRO FRICG_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.3800 0.3200 0.4700 0.5800 ;
        RECT 0.9000 0.3200 0.9900 0.5800 ;
        RECT 1.8000 0.3200 1.9700 0.3900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 1.0950 2.5950 1.1950 ;
        RECT 2.2100 1.0500 2.3900 1.0950 ;
    END
    ANTENNAGATEAREA 0.132 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3200 1.4500 0.9500 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8200 ;
        RECT 0.8600 1.5500 0.9500 1.8200 ;
        RECT 0.3200 0.9300 0.4100 1.4500 ;
        RECT 0.1200 0.8400 0.7300 0.9300 ;
        RECT 0.6400 0.4850 0.7300 0.8400 ;
        RECT 0.1200 0.4700 0.2100 0.8400 ;
    END
    ANTENNADIFFAREA 0.5958 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.0800 1.8400 0.1700 2.0800 ;
        RECT 0.6000 1.8400 0.6900 2.0800 ;
        RECT 1.1200 1.8400 1.2100 2.0800 ;
        RECT 2.3700 1.5250 2.4600 2.0800 ;
        RECT 1.7150 1.2950 1.8050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.2050 0.7100 1.4300 0.8000 ;
      RECT 1.3400 0.4100 1.4300 0.7100 ;
      RECT 1.2700 1.1600 1.9200 1.1950 ;
      RECT 1.1500 1.1050 1.9200 1.1600 ;
      RECT 1.3900 1.1950 1.4800 1.4550 ;
      RECT 1.1500 1.0700 1.3600 1.1050 ;
      RECT 2.0100 1.2850 2.7200 1.3750 ;
      RECT 2.6300 1.3750 2.7200 1.6950 ;
      RECT 0.9500 0.8900 2.5000 0.9600 ;
      RECT 2.0100 0.8700 2.5000 0.8900 ;
      RECT 2.3300 0.6600 2.5000 0.8700 ;
      RECT 0.9500 0.9800 1.0400 1.0900 ;
      RECT 0.5000 1.0900 1.0400 1.1800 ;
      RECT 2.1100 1.4000 2.2000 1.6800 ;
      RECT 2.0100 1.3750 2.2000 1.4000 ;
      RECT 2.0100 0.9800 2.1000 1.2850 ;
      RECT 0.9500 0.9600 2.1000 0.9800 ;
      RECT 1.5700 0.5700 1.6600 0.7800 ;
      RECT 1.5700 0.4800 2.7200 0.5700 ;
      RECT 2.1100 0.5700 2.2000 0.7800 ;
      RECT 2.6300 0.5700 2.7200 0.8500 ;
      RECT 1.5700 0.4100 1.6600 0.4800 ;
      RECT 2.1100 0.4100 2.2000 0.4800 ;
  END
END FRICG_X4B_A12TH

MACRO FRICG_X5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.5950 0.3200 0.6850 0.5700 ;
        RECT 1.1150 0.3200 1.2050 0.5700 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4100 1.2500 2.8300 1.3500 ;
    END
    ANTENNAGATEAREA 0.162 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4500 1.2100 1.5500 ;
        RECT 0.0800 1.5500 0.1700 1.8200 ;
        RECT 0.6000 1.5500 0.6900 1.8200 ;
        RECT 1.1200 1.5500 1.2100 1.8200 ;
        RECT 0.0800 1.0000 0.1700 1.4500 ;
        RECT 0.0800 0.9100 0.9450 1.0000 ;
        RECT 0.3350 0.6100 0.4250 0.9100 ;
        RECT 0.8550 0.6100 0.9450 0.9100 ;
    END
    ANTENNADIFFAREA 0.8022 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.3400 1.8400 0.4300 2.0800 ;
        RECT 0.8600 1.8400 0.9500 2.0800 ;
        RECT 1.3800 1.8400 1.4700 2.0800 ;
        RECT 2.5700 1.8050 2.6600 2.0800 ;
        RECT 1.9600 1.4700 2.0500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.4650 0.6000 1.5550 0.8300 ;
      RECT 1.4650 0.5100 1.6300 0.6000 ;
      RECT 1.5400 0.4100 1.6300 0.5100 ;
      RECT 1.4600 1.1000 2.1000 1.1900 ;
      RECT 1.7000 1.2300 1.7900 1.6550 ;
      RECT 1.4600 1.1900 1.7900 1.2300 ;
      RECT 2.2100 1.4400 2.9200 1.5300 ;
      RECT 2.8300 1.5300 2.9200 1.8500 ;
      RECT 1.1950 0.9200 2.6600 1.0100 ;
      RECT 2.5700 0.6800 2.6600 0.9200 ;
      RECT 1.1950 1.0100 1.2850 1.0900 ;
      RECT 0.4150 1.0900 1.2850 1.1800 ;
      RECT 2.3100 1.5550 2.4000 1.8550 ;
      RECT 2.2100 1.5300 2.4000 1.5550 ;
      RECT 2.2100 1.0100 2.3000 1.4400 ;
      RECT 1.7900 0.5700 1.8800 0.6750 ;
      RECT 1.7900 0.4800 2.9200 0.5700 ;
      RECT 2.3100 0.5700 2.4000 0.8300 ;
      RECT 2.8300 0.5700 2.9200 0.8500 ;
      RECT 2.3100 0.4600 2.4000 0.4800 ;
  END
END FRICG_X5B_A12TH

MACRO FRICG_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9800 ;
        RECT 1.4600 0.3200 1.5500 0.7050 ;
        RECT 1.8250 0.3200 1.9150 0.9150 ;
        RECT 2.3450 0.3200 2.4350 0.7150 ;
        RECT 2.8650 0.3200 2.9550 0.7150 ;
        RECT 3.3850 0.3200 3.4750 0.9350 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 1.0450 1.2050 1.2350 ;
    END
    ANTENNAGATEAREA 0.192 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9500 3.1500 1.2500 ;
        RECT 2.0800 1.2500 3.2150 1.3500 ;
        RECT 2.0850 0.8500 3.2150 0.9500 ;
        RECT 2.0800 1.3500 2.1800 1.7200 ;
        RECT 2.6050 1.3500 2.6950 1.7200 ;
        RECT 3.1250 1.3500 3.2150 1.7000 ;
        RECT 2.6050 0.5700 2.6950 0.8500 ;
        RECT 3.1250 0.5700 3.2150 0.8500 ;
        RECT 2.0850 0.5500 2.1750 0.8500 ;
    END
    ANTENNADIFFAREA 0.876 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 0.7200 1.7700 0.8100 2.0800 ;
        RECT 1.2400 1.7700 1.3300 2.0800 ;
        RECT 1.8250 1.7700 1.9150 2.0800 ;
        RECT 2.3450 1.7700 2.4350 2.0800 ;
        RECT 2.8650 1.7700 2.9550 2.0800 ;
        RECT 3.3850 1.7700 3.4750 2.0800 ;
        RECT 0.0800 1.5800 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7700 0.1700 1.4700 ;
      RECT 0.3400 1.3300 1.4450 1.4200 ;
      RECT 1.3550 1.1750 1.4450 1.3300 ;
      RECT 0.3400 1.4200 0.4300 1.7800 ;
      RECT 0.4800 1.0850 0.5700 1.3300 ;
      RECT 1.6250 1.0550 2.9000 1.1450 ;
      RECT 0.9800 1.6300 1.0700 1.9600 ;
      RECT 0.9300 0.4700 1.0200 0.8100 ;
      RECT 0.9800 1.5400 1.7150 1.6300 ;
      RECT 1.6250 1.1450 1.7150 1.5400 ;
      RECT 1.6250 0.9000 1.7150 1.0550 ;
      RECT 0.9300 0.8100 1.7150 0.9000 ;
  END
END FRICG_X6B_A12TH

MACRO FRICG_X7P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9550 ;
        RECT 1.3750 0.3200 1.4650 0.6950 ;
        RECT 2.1950 0.3200 2.2850 0.6750 ;
        RECT 2.7300 0.3200 2.8200 0.6450 ;
        RECT 3.2500 0.3200 3.3400 0.6450 ;
        RECT 3.7700 0.3200 3.8600 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.6750 1.9500 0.7650 2.0800 ;
        RECT 1.9050 1.7700 1.9950 2.0800 ;
        RECT 2.4700 1.7700 2.5600 2.0800 ;
        RECT 2.9900 1.7700 3.0800 2.0800 ;
        RECT 3.5100 1.7700 3.6000 2.0800 ;
        RECT 1.1950 1.7650 1.2850 2.0800 ;
        RECT 0.0800 1.5400 0.1700 2.0800 ;
    END
  END VDD

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4450 0.8450 3.5550 1.2650 ;
        RECT 2.1700 1.2650 3.8650 1.3750 ;
        RECT 2.4650 0.7350 3.6050 0.8450 ;
        RECT 2.1700 1.3750 2.2700 1.7450 ;
        RECT 2.7250 1.3750 2.8250 1.7450 ;
        RECT 3.2450 1.3750 3.3450 1.7450 ;
        RECT 3.7650 1.3750 3.8650 1.7450 ;
        RECT 2.4650 0.4250 2.5650 0.7350 ;
        RECT 2.9850 0.4250 3.0850 0.7350 ;
        RECT 3.5050 0.4250 3.6050 0.7350 ;
    END
    ANTENNADIFFAREA 1.1615 ;
  END ECK

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.0500 1.8200 1.1500 ;
        RECT 1.7300 1.1500 1.8200 1.2900 ;
    END
    ANTENNAGATEAREA 0.24 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7450 0.1700 1.4300 ;
      RECT 0.3400 1.2500 1.6200 1.3400 ;
      RECT 0.3400 1.3400 0.4300 1.7150 ;
      RECT 0.4450 1.0850 0.5350 1.2500 ;
      RECT 1.9100 0.9600 3.2750 1.0500 ;
      RECT 0.9350 1.6400 1.0250 1.9600 ;
      RECT 0.8300 0.4950 0.9200 0.8500 ;
      RECT 0.9350 1.5500 2.0000 1.6400 ;
      RECT 1.9100 1.0500 2.0000 1.5500 ;
      RECT 1.9100 0.9400 2.0000 0.9600 ;
      RECT 0.8300 0.8500 2.0000 0.9400 ;
      RECT 1.8350 0.5100 1.9250 0.8500 ;
  END
END FRICG_X7P5B_A12TH

MACRO FRICG_X9B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3400 0.3200 0.4300 0.9100 ;
        RECT 1.3750 0.3200 1.4650 0.6300 ;
        RECT 2.1950 0.3200 2.2850 0.6300 ;
        RECT 2.7300 0.3200 2.8200 0.6200 ;
        RECT 3.2500 0.3200 3.3400 0.6200 ;
        RECT 3.7700 0.3200 3.8600 0.6200 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.1000 1.1500 1.1900 ;
        RECT 0.7500 1.0450 1.8200 1.1000 ;
        RECT 1.7300 1.1000 1.8200 1.2850 ;
        RECT 1.0500 1.0000 1.8200 1.0450 ;
    END
    ANTENNAGATEAREA 0.2826 ;
  END CK

  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8350 0.8400 3.9650 1.2350 ;
        RECT 2.1700 1.2350 3.9650 1.3650 ;
        RECT 2.4650 0.7100 4.1250 0.8400 ;
        RECT 2.1700 1.3650 2.2700 1.7150 ;
        RECT 2.7000 1.3650 2.8000 1.7150 ;
        RECT 3.2200 1.3650 3.3200 1.7150 ;
        RECT 3.7400 1.3650 3.8400 1.7150 ;
        RECT 2.4650 0.4200 2.5650 0.7100 ;
        RECT 2.9850 0.4200 3.0850 0.7100 ;
        RECT 3.5050 0.4200 3.6050 0.7100 ;
        RECT 4.0250 0.4200 4.1250 0.7100 ;
    END
    ANTENNADIFFAREA 1.32355 ;
  END ECK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.6750 1.9650 0.7650 2.0800 ;
        RECT 1.9050 1.7700 1.9950 2.0800 ;
        RECT 2.4450 1.7700 2.5350 2.0800 ;
        RECT 2.9650 1.7700 3.0550 2.0800 ;
        RECT 3.4850 1.7700 3.5750 2.0800 ;
        RECT 4.0300 1.7700 4.1200 2.0800 ;
        RECT 1.1950 1.7450 1.2850 2.0800 ;
        RECT 0.0800 1.6650 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 0.7000 0.1700 1.5150 ;
      RECT 0.3400 1.3300 1.3300 1.4200 ;
      RECT 1.2400 1.3000 1.3300 1.3300 ;
      RECT 1.2400 1.2100 1.6300 1.3000 ;
      RECT 0.3400 1.4200 0.4300 1.7750 ;
      RECT 0.4800 1.0850 0.5700 1.3300 ;
      RECT 1.9100 0.9300 3.6050 1.0200 ;
      RECT 0.9350 1.6400 1.0250 1.9600 ;
      RECT 0.8450 0.4700 0.9350 0.8100 ;
      RECT 0.9350 1.5500 2.0000 1.6400 ;
      RECT 1.9100 1.0200 2.0000 1.5500 ;
      RECT 1.9100 0.9000 2.0000 0.9300 ;
      RECT 0.8450 0.8100 2.0000 0.9000 ;
      RECT 1.8350 0.4150 1.9250 0.8100 ;
  END
END FRICG_X9B_A12TH

MACRO FILL64_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.8450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.8450 0.3200 ;
    END
  END VSS
END FILL64_A12TH

MACRO FILL8_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
    END
  END VSS
END FILL8_A12TH

MACRO FILLCAP128_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 25.6450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
        RECT 2.6900 1.7700 2.7900 2.0800 ;
        RECT 3.2100 1.7700 3.3100 2.0800 ;
        RECT 3.7300 1.7700 3.8300 2.0800 ;
        RECT 4.2500 1.7700 4.3500 2.0800 ;
        RECT 4.7700 1.7700 4.8700 2.0800 ;
        RECT 5.2900 1.7700 5.3900 2.0800 ;
        RECT 5.8100 1.7700 5.9100 2.0800 ;
        RECT 6.8500 1.7700 6.9500 2.0800 ;
        RECT 7.3700 1.7700 7.4700 2.0800 ;
        RECT 7.8900 1.7700 7.9900 2.0800 ;
        RECT 8.4100 1.7700 8.5100 2.0800 ;
        RECT 6.3300 1.7550 6.4300 2.0800 ;
        RECT 8.9300 1.7700 9.0300 2.0800 ;
        RECT 9.4500 1.7700 9.5500 2.0800 ;
        RECT 9.9700 1.7700 10.0700 2.0800 ;
        RECT 10.4900 1.7700 10.5900 2.0800 ;
        RECT 11.0100 1.7700 11.1100 2.0800 ;
        RECT 11.5300 1.7700 11.6300 2.0800 ;
        RECT 12.0500 1.7700 12.1500 2.0800 ;
        RECT 12.5700 1.7700 12.6700 2.0800 ;
        RECT 13.0900 1.7700 13.1900 2.0800 ;
        RECT 13.6100 1.7700 13.7100 2.0800 ;
        RECT 14.1300 1.7700 14.2300 2.0800 ;
        RECT 14.6500 1.7700 14.7500 2.0800 ;
        RECT 15.1700 1.7700 15.2700 2.0800 ;
        RECT 15.6900 1.7700 15.7900 2.0800 ;
        RECT 16.2100 1.7700 16.3100 2.0800 ;
        RECT 16.7300 1.7700 16.8300 2.0800 ;
        RECT 17.2500 1.7700 17.3500 2.0800 ;
        RECT 17.7700 1.7700 17.8700 2.0800 ;
        RECT 18.2900 1.7700 18.3900 2.0800 ;
        RECT 19.3300 1.7700 19.4300 2.0800 ;
        RECT 19.8500 1.7700 19.9500 2.0800 ;
        RECT 20.3700 1.7700 20.4700 2.0800 ;
        RECT 20.8900 1.7700 20.9900 2.0800 ;
        RECT 21.4100 1.7700 21.5100 2.0800 ;
        RECT 21.9300 1.7700 22.0300 2.0800 ;
        RECT 22.4500 1.7700 22.5500 2.0800 ;
        RECT 22.9700 1.7700 23.0700 2.0800 ;
        RECT 23.4900 1.7700 23.5900 2.0800 ;
        RECT 24.0100 1.7700 24.1100 2.0800 ;
        RECT 24.5300 1.7700 24.6300 2.0800 ;
        RECT 25.0500 1.7700 25.1500 2.0800 ;
        RECT 18.8100 1.7550 18.9100 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 25.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6600 ;
        RECT 0.6100 0.3200 0.7100 0.6600 ;
        RECT 1.1300 0.3200 1.2300 0.6600 ;
        RECT 1.6500 0.3200 1.7500 0.6600 ;
        RECT 2.1700 0.3200 2.2700 0.6600 ;
        RECT 2.6900 0.3200 2.7900 0.6600 ;
        RECT 3.2100 0.3200 3.3100 0.6600 ;
        RECT 3.7300 0.3200 3.8300 0.6600 ;
        RECT 4.2500 0.3200 4.3500 0.6600 ;
        RECT 4.7700 0.3200 4.8700 0.6600 ;
        RECT 5.2900 0.3200 5.3900 0.6600 ;
        RECT 5.8100 0.3200 5.9100 0.6600 ;
        RECT 6.3300 0.3200 6.4300 0.6600 ;
        RECT 6.8500 0.3200 6.9500 0.6600 ;
        RECT 7.3700 0.3200 7.4700 0.6600 ;
        RECT 7.8900 0.3200 7.9900 0.6600 ;
        RECT 8.4100 0.3200 8.5100 0.6600 ;
        RECT 8.9300 0.3200 9.0300 0.6600 ;
        RECT 9.4500 0.3200 9.5500 0.6600 ;
        RECT 9.9700 0.3200 10.0700 0.6600 ;
        RECT 10.4900 0.3200 10.5900 0.6600 ;
        RECT 11.0100 0.3200 11.1100 0.6600 ;
        RECT 11.5300 0.3200 11.6300 0.6600 ;
        RECT 12.0500 0.3200 12.1500 0.6600 ;
        RECT 12.5700 0.3200 12.6700 0.6600 ;
        RECT 13.0900 0.3200 13.1900 0.6600 ;
        RECT 13.6100 0.3200 13.7100 0.6600 ;
        RECT 14.1300 0.3200 14.2300 0.6600 ;
        RECT 14.6500 0.3200 14.7500 0.6600 ;
        RECT 15.1700 0.3200 15.2700 0.6600 ;
        RECT 15.6900 0.3200 15.7900 0.6600 ;
        RECT 16.2100 0.3200 16.3100 0.6600 ;
        RECT 16.7300 0.3200 16.8300 0.6600 ;
        RECT 17.2500 0.3200 17.3500 0.6600 ;
        RECT 17.7700 0.3200 17.8700 0.6600 ;
        RECT 18.2900 0.3200 18.3900 0.6600 ;
        RECT 18.8100 0.3200 18.9100 0.6600 ;
        RECT 19.3300 0.3200 19.4300 0.6600 ;
        RECT 19.8500 0.3200 19.9500 0.6600 ;
        RECT 20.3700 0.3200 20.4700 0.6600 ;
        RECT 20.8900 0.3200 20.9900 0.6600 ;
        RECT 21.4100 0.3200 21.5100 0.6600 ;
        RECT 21.9300 0.3200 22.0300 0.6600 ;
        RECT 22.4500 0.3200 22.5500 0.6600 ;
        RECT 22.9700 0.3200 23.0700 0.6600 ;
        RECT 23.4900 0.3200 23.5900 0.6600 ;
        RECT 24.0100 0.3200 24.1100 0.6600 ;
        RECT 24.5300 0.3200 24.6300 0.6600 ;
        RECT 25.0500 0.3200 25.1500 0.6600 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.4750 25.4050 1.5650 ;
      RECT 25.3150 1.5650 25.4050 1.9050 ;
      RECT 0.3550 1.0050 25.0600 1.0950 ;
      RECT 0.3550 1.0950 0.4450 1.4750 ;
      RECT 0.3550 1.5650 0.4450 1.9050 ;
      RECT 0.8750 1.5650 0.9650 1.9050 ;
      RECT 1.3950 1.5650 1.4850 1.9050 ;
      RECT 1.9150 1.5650 2.0050 1.9050 ;
      RECT 2.4350 1.5650 2.5250 1.9050 ;
      RECT 2.9550 1.5650 3.0450 1.9050 ;
      RECT 3.4750 1.5650 3.5650 1.9050 ;
      RECT 3.9950 1.5650 4.0850 1.9050 ;
      RECT 4.5150 1.5650 4.6050 1.9050 ;
      RECT 5.0350 1.5650 5.1250 1.9050 ;
      RECT 5.5550 1.5650 5.6450 1.9050 ;
      RECT 6.0750 1.5650 6.1650 1.9050 ;
      RECT 6.5950 1.5650 6.6850 1.9050 ;
      RECT 7.1150 1.5650 7.2050 1.9050 ;
      RECT 7.6350 1.5650 7.7250 1.9050 ;
      RECT 8.1550 1.5650 8.2450 1.9050 ;
      RECT 8.6750 1.5650 8.7650 1.9050 ;
      RECT 9.1950 1.5650 9.2850 1.9050 ;
      RECT 9.7150 1.5650 9.8050 1.9050 ;
      RECT 10.2350 1.5650 10.3250 1.9050 ;
      RECT 10.7550 1.5650 10.8450 1.9050 ;
      RECT 11.2750 1.5650 11.3650 1.9050 ;
      RECT 11.7950 1.5650 11.8850 1.9050 ;
      RECT 12.3150 1.5650 12.4050 1.9050 ;
      RECT 12.8350 1.5650 12.9250 1.9300 ;
      RECT 13.3550 1.5650 13.4450 1.9050 ;
      RECT 13.8750 1.5650 13.9650 1.9050 ;
      RECT 14.3950 1.5650 14.4850 1.9050 ;
      RECT 14.9150 1.5650 15.0050 1.9050 ;
      RECT 15.4350 1.5650 15.5250 1.9050 ;
      RECT 15.9550 1.5650 16.0450 1.9050 ;
      RECT 16.4750 1.5650 16.5650 1.9050 ;
      RECT 16.9950 1.5650 17.0850 1.9050 ;
      RECT 17.5150 1.5650 17.6050 1.9050 ;
      RECT 18.0350 1.5650 18.1250 1.9050 ;
      RECT 18.5550 1.5650 18.6450 1.9050 ;
      RECT 19.0750 1.5650 19.1650 1.9050 ;
      RECT 19.5950 1.5650 19.6850 1.9050 ;
      RECT 20.1150 1.5650 20.2050 1.9050 ;
      RECT 20.6350 1.5650 20.7250 1.9050 ;
      RECT 21.1550 1.5650 21.2450 1.9050 ;
      RECT 21.6750 1.5650 21.7650 1.9050 ;
      RECT 22.1950 1.5650 22.2850 1.9050 ;
      RECT 22.7150 1.5650 22.8050 1.9050 ;
      RECT 23.2350 1.5650 23.3250 1.9050 ;
      RECT 23.7550 1.5650 23.8450 1.9050 ;
      RECT 24.2750 1.5650 24.3650 1.9050 ;
      RECT 24.7950 1.5650 24.8850 1.9050 ;
      RECT 0.6700 1.2650 25.4050 1.3550 ;
      RECT 25.3150 0.8850 25.4050 1.2650 ;
      RECT 0.3550 0.7950 25.4050 0.8850 ;
      RECT 25.3150 0.4550 25.4050 0.7950 ;
      RECT 0.3550 0.4550 0.4450 0.7950 ;
      RECT 0.8750 0.4550 0.9650 0.7950 ;
      RECT 1.3950 0.4550 1.4850 0.7950 ;
      RECT 1.9150 0.4550 2.0050 0.7950 ;
      RECT 2.4350 0.4550 2.5250 0.7950 ;
      RECT 2.9550 0.4550 3.0450 0.7950 ;
      RECT 3.4750 0.4550 3.5650 0.7950 ;
      RECT 3.9950 0.4550 4.0850 0.7950 ;
      RECT 4.5150 0.4550 4.6050 0.7950 ;
      RECT 5.0350 0.4550 5.1250 0.7950 ;
      RECT 5.5550 0.4550 5.6450 0.7950 ;
      RECT 6.0750 0.4550 6.1650 0.7950 ;
      RECT 6.5950 0.4550 6.6850 0.7950 ;
      RECT 7.1150 0.4550 7.2050 0.7950 ;
      RECT 7.6350 0.4550 7.7250 0.7950 ;
      RECT 8.1550 0.4550 8.2450 0.7950 ;
      RECT 8.6750 0.4550 8.7650 0.7950 ;
      RECT 9.1950 0.4550 9.2850 0.7950 ;
      RECT 9.7150 0.4550 9.8050 0.7950 ;
      RECT 10.2350 0.4550 10.3250 0.7950 ;
      RECT 10.7550 0.4550 10.8450 0.7950 ;
      RECT 11.2750 0.4550 11.3650 0.7950 ;
      RECT 11.7950 0.4550 11.8850 0.7950 ;
      RECT 12.3150 0.4550 12.4050 0.7950 ;
      RECT 12.8350 0.4550 12.9250 0.7950 ;
      RECT 13.3550 0.4550 13.4450 0.7950 ;
      RECT 13.8750 0.4550 13.9650 0.7950 ;
      RECT 14.3950 0.4550 14.4850 0.7950 ;
      RECT 14.9150 0.4550 15.0050 0.7950 ;
      RECT 15.4350 0.4550 15.5250 0.7950 ;
      RECT 15.9550 0.4550 16.0450 0.7950 ;
      RECT 16.4750 0.4550 16.5650 0.7950 ;
      RECT 16.9950 0.4550 17.0850 0.7950 ;
      RECT 17.5150 0.4550 17.6050 0.7950 ;
      RECT 18.0350 0.4550 18.1250 0.7950 ;
      RECT 18.5550 0.4550 18.6450 0.7950 ;
      RECT 19.0750 0.4550 19.1650 0.7950 ;
      RECT 19.5950 0.4550 19.6850 0.7950 ;
      RECT 20.1150 0.4550 20.2050 0.7950 ;
      RECT 20.6350 0.4550 20.7250 0.7950 ;
      RECT 21.1550 0.4550 21.2450 0.7950 ;
      RECT 21.6750 0.4550 21.7650 0.7950 ;
      RECT 22.1950 0.4550 22.2850 0.7950 ;
      RECT 22.7150 0.4550 22.8050 0.7950 ;
      RECT 23.2350 0.4550 23.3250 0.7950 ;
      RECT 23.7550 0.4550 23.8450 0.7950 ;
      RECT 24.2750 0.4550 24.3650 0.7950 ;
      RECT 24.7950 0.4550 24.8850 0.7950 ;
  END
END FILLCAP128_A12TH

MACRO FILLCAP16_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
        RECT 2.6900 1.7700 2.7900 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
        RECT 1.1300 0.3200 1.2300 0.6300 ;
        RECT 1.6500 0.3200 1.7500 0.6300 ;
        RECT 2.1700 0.3200 2.2700 0.6300 ;
        RECT 2.6900 0.3200 2.7900 0.6300 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.4750 3.0450 1.5650 ;
      RECT 2.9550 1.5650 3.0450 1.9050 ;
      RECT 0.3550 1.5650 0.4450 1.9050 ;
      RECT 0.3550 1.0950 0.4450 1.4750 ;
      RECT 0.8750 1.5650 0.9650 1.9050 ;
      RECT 1.3950 1.5650 1.4850 1.9050 ;
      RECT 1.9150 1.5650 2.0050 1.9050 ;
      RECT 2.4350 1.5650 2.5250 1.9050 ;
      RECT 0.3550 1.0050 2.4400 1.0950 ;
      RECT 0.6700 1.2650 2.6950 1.3550 ;
      RECT 2.6050 0.8850 2.6950 1.2650 ;
      RECT 0.3550 0.7950 3.0450 0.8850 ;
      RECT 2.9550 0.4550 3.0450 0.7950 ;
      RECT 0.3550 0.4550 0.4450 0.7950 ;
      RECT 0.8750 0.4550 0.9650 0.7950 ;
      RECT 1.3950 0.4550 1.4850 0.7950 ;
      RECT 1.9150 0.4550 2.0050 0.7950 ;
      RECT 2.4350 0.4550 2.5250 0.7950 ;
  END
END FILLCAP16_A12TH

MACRO FILLCAP32_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
        RECT 2.6900 1.7700 2.7900 2.0800 ;
        RECT 3.2100 1.7700 3.3100 2.0800 ;
        RECT 3.7300 1.7700 3.8300 2.0800 ;
        RECT 4.2500 1.7700 4.3500 2.0800 ;
        RECT 4.7700 1.7700 4.8700 2.0800 ;
        RECT 5.2900 1.7700 5.3900 2.0800 ;
        RECT 5.8100 1.7700 5.9100 2.0800 ;
        RECT 6.3300 1.7700 6.4300 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
        RECT 1.1300 0.3200 1.2300 0.6300 ;
        RECT 1.6500 0.3200 1.7500 0.6300 ;
        RECT 2.1700 0.3200 2.2700 0.6300 ;
        RECT 2.6900 0.3200 2.7900 0.6300 ;
        RECT 3.2100 0.3200 3.3100 0.6300 ;
        RECT 3.7300 0.3200 3.8300 0.6300 ;
        RECT 4.2500 0.3200 4.3500 0.6300 ;
        RECT 4.7700 0.3200 4.8700 0.6300 ;
        RECT 5.2900 0.3200 5.3900 0.6300 ;
        RECT 5.8100 0.3200 5.9100 0.6300 ;
        RECT 6.3300 0.3200 6.4300 0.6300 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.4750 6.1650 1.5650 ;
      RECT 6.0750 1.5650 6.1650 1.9050 ;
      RECT 0.3550 1.5650 0.4450 1.9050 ;
      RECT 0.3550 1.0950 0.4450 1.4750 ;
      RECT 0.8750 1.5650 0.9650 1.9050 ;
      RECT 1.3950 1.5650 1.4850 1.9050 ;
      RECT 1.9150 1.5650 2.0050 1.9050 ;
      RECT 2.4350 1.5650 2.5250 1.9050 ;
      RECT 2.9550 1.5650 3.0450 1.9050 ;
      RECT 3.4750 1.5650 3.5650 1.9050 ;
      RECT 3.9950 1.5650 4.0850 1.9050 ;
      RECT 4.5150 1.5650 4.6050 1.9050 ;
      RECT 5.0350 1.5650 5.1250 1.9050 ;
      RECT 5.5550 1.5650 5.6450 1.9050 ;
      RECT 0.3550 1.0050 5.5600 1.0950 ;
      RECT 0.6700 1.2650 6.1650 1.3550 ;
      RECT 6.0750 0.8850 6.1650 1.2650 ;
      RECT 0.3550 0.7950 6.1650 0.8850 ;
      RECT 6.0750 0.4550 6.1650 0.7950 ;
      RECT 0.3550 0.4550 0.4450 0.7950 ;
      RECT 0.8750 0.4550 0.9650 0.7950 ;
      RECT 1.3950 0.4550 1.4850 0.7950 ;
      RECT 1.9150 0.4550 2.0050 0.7950 ;
      RECT 2.4350 0.4550 2.5250 0.7950 ;
      RECT 2.9550 0.4550 3.0450 0.7950 ;
      RECT 3.4750 0.4550 3.5650 0.7950 ;
      RECT 3.9950 0.4550 4.0850 0.7950 ;
      RECT 4.5150 0.4550 4.6050 0.7950 ;
      RECT 5.0350 0.4550 5.1250 0.7950 ;
      RECT 5.5550 0.4550 5.6450 0.7950 ;
  END
END FILLCAP32_A12TH

MACRO FILLCAP3_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.6450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.6450 0.3200 ;
        RECT 0.1000 0.3200 0.2000 0.6300 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0950 1.0400 0.1850 1.8400 ;
      RECT 0.0950 0.9500 0.2750 1.0400 ;
      RECT 0.3650 0.4100 0.4550 1.3600 ;
  END
END FILLCAP3_A12TH

MACRO FILLCAP4_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.5100 0.4450 1.8500 ;
      RECT 0.2150 1.4200 0.4450 1.5100 ;
      RECT 0.2150 1.0400 0.3050 1.4200 ;
      RECT 0.0750 0.9500 0.3050 1.0400 ;
      RECT 0.4250 1.2100 0.6950 1.3000 ;
      RECT 0.4250 0.8400 0.5150 1.2100 ;
      RECT 0.3550 0.7500 0.5150 0.8400 ;
      RECT 0.3550 0.4100 0.4450 0.7500 ;
  END
END FILLCAP4_A12TH

MACRO FILLCAP64_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.8450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
        RECT 2.6900 1.7700 2.7900 2.0800 ;
        RECT 3.2100 1.7700 3.3100 2.0800 ;
        RECT 3.7300 1.7700 3.8300 2.0800 ;
        RECT 4.2500 1.7700 4.3500 2.0800 ;
        RECT 4.7700 1.7700 4.8700 2.0800 ;
        RECT 5.2900 1.7700 5.3900 2.0800 ;
        RECT 5.8100 1.7700 5.9100 2.0800 ;
        RECT 6.3300 1.7700 6.4300 2.0800 ;
        RECT 6.8500 1.7700 6.9500 2.0800 ;
        RECT 7.3700 1.7700 7.4700 2.0800 ;
        RECT 7.8900 1.7700 7.9900 2.0800 ;
        RECT 8.4100 1.7700 8.5100 2.0800 ;
        RECT 8.9300 1.7700 9.0300 2.0800 ;
        RECT 9.4500 1.7700 9.5500 2.0800 ;
        RECT 9.9700 1.7700 10.0700 2.0800 ;
        RECT 10.4900 1.7700 10.5900 2.0800 ;
        RECT 11.0100 1.7700 11.1100 2.0800 ;
        RECT 11.5300 1.7700 11.6300 2.0800 ;
        RECT 12.0500 1.7700 12.1500 2.0800 ;
        RECT 12.5700 1.7700 12.6700 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6800 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
        RECT 1.1300 0.3200 1.2300 0.6300 ;
        RECT 1.6500 0.3200 1.7500 0.6300 ;
        RECT 2.1700 0.3200 2.2700 0.6300 ;
        RECT 2.6900 0.3200 2.7900 0.6300 ;
        RECT 3.2100 0.3200 3.3100 0.6300 ;
        RECT 3.7300 0.3200 3.8300 0.6300 ;
        RECT 4.2500 0.3200 4.3500 0.6300 ;
        RECT 4.7700 0.3200 4.8700 0.6300 ;
        RECT 5.2900 0.3200 5.3900 0.6300 ;
        RECT 5.8100 0.3200 5.9100 0.6300 ;
        RECT 6.3300 0.3200 6.4300 0.6300 ;
        RECT 6.8500 0.3200 6.9500 0.6300 ;
        RECT 7.3700 0.3200 7.4700 0.6300 ;
        RECT 7.8900 0.3200 7.9900 0.6300 ;
        RECT 8.4100 0.3200 8.5100 0.6300 ;
        RECT 8.9300 0.3200 9.0300 0.6300 ;
        RECT 9.4500 0.3200 9.5500 0.6300 ;
        RECT 9.9700 0.3200 10.0700 0.6300 ;
        RECT 10.4900 0.3200 10.5900 0.6300 ;
        RECT 11.0100 0.3200 11.1100 0.6300 ;
        RECT 11.5300 0.3200 11.6300 0.6300 ;
        RECT 12.0500 0.3200 12.1500 0.6300 ;
        RECT 12.5700 0.3200 12.6700 0.6300 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.4750 12.4050 1.5650 ;
      RECT 12.3150 1.5650 12.4050 1.9050 ;
      RECT 0.3550 1.5650 0.4450 1.9050 ;
      RECT 0.3550 1.0950 0.4450 1.4750 ;
      RECT 0.8750 1.5650 0.9650 1.9050 ;
      RECT 1.3950 1.5650 1.4850 1.9050 ;
      RECT 1.9150 1.5650 2.0050 1.9050 ;
      RECT 2.4350 1.5650 2.5250 1.9050 ;
      RECT 2.9550 1.5650 3.0450 1.9050 ;
      RECT 3.4750 1.5650 3.5650 1.9050 ;
      RECT 3.9950 1.5650 4.0850 1.9050 ;
      RECT 4.5150 1.5650 4.6050 1.9050 ;
      RECT 5.0350 1.5650 5.1250 1.9050 ;
      RECT 5.5550 1.5650 5.6450 1.9050 ;
      RECT 6.0750 1.5650 6.1650 1.9050 ;
      RECT 6.5950 1.5650 6.6850 1.9050 ;
      RECT 7.1150 1.5650 7.2050 1.9050 ;
      RECT 7.6350 1.5650 7.7250 1.9050 ;
      RECT 8.1550 1.5650 8.2450 1.9050 ;
      RECT 8.6750 1.5650 8.7650 1.9050 ;
      RECT 9.1950 1.5650 9.2850 1.9050 ;
      RECT 9.7150 1.5650 9.8050 1.9050 ;
      RECT 10.2350 1.5650 10.3250 1.9050 ;
      RECT 10.7550 1.5650 10.8450 1.9050 ;
      RECT 11.2750 1.5650 11.3650 1.9050 ;
      RECT 11.7950 1.5650 11.8850 1.9050 ;
      RECT 0.3550 1.0050 11.8000 1.0950 ;
      RECT 0.6700 1.2650 12.4050 1.3550 ;
      RECT 12.3150 0.8850 12.4050 1.2650 ;
      RECT 0.3550 0.7950 12.4050 0.8850 ;
      RECT 12.3150 0.4550 12.4050 0.7950 ;
      RECT 0.3550 0.4550 0.4450 0.7950 ;
      RECT 0.8750 0.4550 0.9650 0.7950 ;
      RECT 1.3950 0.4550 1.4850 0.7950 ;
      RECT 1.9150 0.4550 2.0050 0.7950 ;
      RECT 2.4350 0.4550 2.5250 0.7950 ;
      RECT 2.9550 0.4550 3.0450 0.7950 ;
      RECT 3.4750 0.4550 3.5650 0.7950 ;
      RECT 3.9950 0.4550 4.0850 0.7950 ;
      RECT 4.5150 0.4550 4.6050 0.7950 ;
      RECT 5.0350 0.4550 5.1250 0.7950 ;
      RECT 5.5550 0.4550 5.6450 0.7950 ;
      RECT 6.0750 0.4550 6.1650 0.7950 ;
      RECT 6.5950 0.4550 6.6850 0.7950 ;
      RECT 7.1150 0.4550 7.2050 0.7950 ;
      RECT 7.6350 0.4550 7.7250 0.7950 ;
      RECT 8.1550 0.4550 8.2450 0.7950 ;
      RECT 8.6750 0.4550 8.7650 0.7950 ;
      RECT 9.1950 0.4550 9.2850 0.7950 ;
      RECT 9.7150 0.4550 9.8050 0.7950 ;
      RECT 10.2350 0.4550 10.3250 0.7950 ;
      RECT 10.7550 0.4550 10.8450 0.7950 ;
      RECT 11.2750 0.4550 11.3650 0.7950 ;
      RECT 11.7950 0.4550 11.8850 0.7950 ;
  END
END FILLCAP64_A12TH

MACRO FILLCAP8_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.0900 1.7550 0.1900 2.0800 ;
        RECT 0.6100 1.7550 0.7100 2.0800 ;
        RECT 1.1300 1.7550 1.2300 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
        RECT 1.1300 0.3200 1.2300 0.6300 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.4750 1.4850 1.5650 ;
      RECT 1.3950 1.5650 1.4850 1.8850 ;
      RECT 0.3550 1.5650 0.4450 1.8850 ;
      RECT 0.3550 1.0950 0.4450 1.4750 ;
      RECT 0.8750 1.5650 0.9650 1.8850 ;
      RECT 0.3550 1.0050 1.0050 1.0950 ;
      RECT 0.5800 1.2650 1.2600 1.3550 ;
      RECT 1.1700 0.8850 1.2600 1.2650 ;
      RECT 0.3550 0.7950 1.4850 0.8850 ;
      RECT 1.3950 0.4750 1.4850 0.7950 ;
      RECT 0.3550 0.4750 0.4450 0.7950 ;
      RECT 0.8750 0.4750 0.9650 0.7950 ;
  END
END FILLCAP8_A12TH

MACRO FILLCAPTIE128_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 25.6450 2.7200 ;
        RECT 0.5100 1.7700 0.6100 2.0800 ;
        RECT 1.0300 1.7700 1.1300 2.0800 ;
        RECT 1.5500 1.7700 1.6500 2.0800 ;
        RECT 0.1350 1.4050 0.2350 2.0800 ;
        RECT 2.0700 1.7700 2.1700 2.0800 ;
        RECT 2.5900 1.7700 2.6900 2.0800 ;
        RECT 3.1100 1.7700 3.2100 2.0800 ;
        RECT 3.6300 1.7700 3.7300 2.0800 ;
        RECT 4.1500 1.7700 4.2500 2.0800 ;
        RECT 4.6700 1.7700 4.7700 2.0800 ;
        RECT 5.1900 1.7700 5.2900 2.0800 ;
        RECT 5.7100 1.7700 5.8100 2.0800 ;
        RECT 6.2300 1.7700 6.3300 2.0800 ;
        RECT 6.7500 1.7700 6.8500 2.0800 ;
        RECT 7.2700 1.7700 7.3700 2.0800 ;
        RECT 7.7900 1.7700 7.8900 2.0800 ;
        RECT 8.3100 1.7700 8.4100 2.0800 ;
        RECT 8.8300 1.7700 8.9300 2.0800 ;
        RECT 9.3500 1.7700 9.4500 2.0800 ;
        RECT 9.8700 1.7700 9.9700 2.0800 ;
        RECT 10.3900 1.7700 10.4900 2.0800 ;
        RECT 10.9100 1.7700 11.0100 2.0800 ;
        RECT 11.4300 1.7700 11.5300 2.0800 ;
        RECT 11.9500 1.7700 12.0500 2.0800 ;
        RECT 12.4700 1.7700 12.5700 2.0800 ;
        RECT 12.9900 1.7700 13.0900 2.0800 ;
        RECT 13.5100 1.7700 13.6100 2.0800 ;
        RECT 14.0300 1.7700 14.1300 2.0800 ;
        RECT 14.5500 1.7700 14.6500 2.0800 ;
        RECT 15.0700 1.7700 15.1700 2.0800 ;
        RECT 15.5900 1.7700 15.6900 2.0800 ;
        RECT 16.1100 1.7700 16.2100 2.0800 ;
        RECT 16.6300 1.7700 16.7300 2.0800 ;
        RECT 17.1500 1.7700 17.2500 2.0800 ;
        RECT 17.6700 1.7700 17.7700 2.0800 ;
        RECT 18.1900 1.7700 18.2900 2.0800 ;
        RECT 18.7100 1.7700 18.8100 2.0800 ;
        RECT 19.2300 1.7700 19.3300 2.0800 ;
        RECT 19.7500 1.7700 19.8500 2.0800 ;
        RECT 20.2700 1.7700 20.3700 2.0800 ;
        RECT 20.7900 1.7700 20.8900 2.0800 ;
        RECT 21.3100 1.7700 21.4100 2.0800 ;
        RECT 21.8300 1.7700 21.9300 2.0800 ;
        RECT 22.3500 1.7700 22.4500 2.0800 ;
        RECT 22.8700 1.7700 22.9700 2.0800 ;
        RECT 23.3900 1.7700 23.4900 2.0800 ;
        RECT 23.9100 1.7700 24.0100 2.0800 ;
        RECT 24.4300 1.7700 24.5300 2.0800 ;
        RECT 24.9500 1.7700 25.0500 2.0800 ;
        RECT 25.3650 1.4050 25.4650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 25.6450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.9750 ;
        RECT 0.5100 0.3200 0.6100 0.6300 ;
        RECT 1.0300 0.3200 1.1300 0.6300 ;
        RECT 1.5500 0.3200 1.6500 0.6300 ;
        RECT 2.0700 0.3200 2.1700 0.6300 ;
        RECT 2.5900 0.3200 2.6900 0.6300 ;
        RECT 3.1100 0.3200 3.2100 0.6300 ;
        RECT 3.6300 0.3200 3.7300 0.6300 ;
        RECT 4.1500 0.3200 4.2500 0.6300 ;
        RECT 4.6700 0.3200 4.7700 0.6300 ;
        RECT 5.1900 0.3200 5.2900 0.6300 ;
        RECT 5.7100 0.3200 5.8100 0.6300 ;
        RECT 6.2300 0.3200 6.3300 0.6300 ;
        RECT 6.7500 0.3200 6.8500 0.6300 ;
        RECT 7.2700 0.3200 7.3700 0.6300 ;
        RECT 7.7900 0.3200 7.8900 0.6300 ;
        RECT 8.3100 0.3200 8.4100 0.6300 ;
        RECT 8.8300 0.3200 8.9300 0.6300 ;
        RECT 9.3500 0.3200 9.4500 0.6300 ;
        RECT 9.8700 0.3200 9.9700 0.6300 ;
        RECT 10.3900 0.3200 10.4900 0.6300 ;
        RECT 10.9100 0.3200 11.0100 0.6300 ;
        RECT 11.4300 0.3200 11.5300 0.6300 ;
        RECT 11.9500 0.3200 12.0500 0.6300 ;
        RECT 12.4700 0.3200 12.5700 0.6300 ;
        RECT 12.9900 0.3200 13.0900 0.6300 ;
        RECT 13.5100 0.3200 13.6100 0.6300 ;
        RECT 14.0300 0.3200 14.1300 0.6300 ;
        RECT 14.5500 0.3200 14.6500 0.6300 ;
        RECT 15.0700 0.3200 15.1700 0.6300 ;
        RECT 15.5900 0.3200 15.6900 0.6300 ;
        RECT 16.1100 0.3200 16.2100 0.6300 ;
        RECT 16.6300 0.3200 16.7300 0.6300 ;
        RECT 17.1500 0.3200 17.2500 0.6300 ;
        RECT 17.6700 0.3200 17.7700 0.6300 ;
        RECT 18.1900 0.3200 18.2900 0.6300 ;
        RECT 18.7100 0.3200 18.8100 0.6300 ;
        RECT 19.2300 0.3200 19.3300 0.6300 ;
        RECT 19.7500 0.3200 19.8500 0.6300 ;
        RECT 20.2700 0.3200 20.3700 0.6300 ;
        RECT 20.7900 0.3200 20.8900 0.6300 ;
        RECT 21.3100 0.3200 21.4100 0.6300 ;
        RECT 21.8300 0.3200 21.9300 0.6300 ;
        RECT 22.3500 0.3200 22.4500 0.6300 ;
        RECT 22.8700 0.3200 22.9700 0.6300 ;
        RECT 23.3900 0.3200 23.4900 0.6300 ;
        RECT 23.9100 0.3200 24.0100 0.6300 ;
        RECT 24.4300 0.3200 24.5300 0.6300 ;
        RECT 24.9500 0.3200 25.0500 0.6300 ;
        RECT 25.3650 0.3200 25.4650 0.9750 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.7750 1.4750 24.7850 1.5650 ;
      RECT 24.6950 1.5650 24.7850 1.8850 ;
      RECT 0.7750 1.0050 24.4650 1.0950 ;
      RECT 0.7750 1.0950 0.8650 1.4750 ;
      RECT 0.7750 1.5650 0.8650 1.9050 ;
      RECT 1.2950 1.5650 1.3850 1.9050 ;
      RECT 1.8150 1.5650 1.9050 1.9050 ;
      RECT 2.3350 1.5650 2.4250 1.9050 ;
      RECT 2.8550 1.5650 2.9450 1.9050 ;
      RECT 3.3750 1.5650 3.4650 1.9050 ;
      RECT 3.8950 1.5650 3.9850 1.9050 ;
      RECT 4.4150 1.5650 4.5050 1.9050 ;
      RECT 4.9350 1.5650 5.0250 1.9050 ;
      RECT 5.4550 1.5650 5.5450 1.9050 ;
      RECT 5.9750 1.5650 6.0650 1.9050 ;
      RECT 6.4950 1.5650 6.5850 1.9050 ;
      RECT 7.0150 1.5650 7.1050 1.9050 ;
      RECT 7.5350 1.5650 7.6250 1.9050 ;
      RECT 8.0550 1.5650 8.1450 1.9050 ;
      RECT 8.5750 1.5650 8.6650 1.9050 ;
      RECT 9.0950 1.5650 9.1850 1.9050 ;
      RECT 9.6150 1.5650 9.7050 1.9050 ;
      RECT 10.1350 1.5650 10.2250 1.9050 ;
      RECT 10.6550 1.5650 10.7450 1.9050 ;
      RECT 11.1750 1.5650 11.2650 1.9050 ;
      RECT 11.6950 1.5650 11.7850 1.9050 ;
      RECT 12.2150 1.5650 12.3050 1.9050 ;
      RECT 12.7350 1.5650 12.8250 1.9050 ;
      RECT 13.2550 1.5650 13.3450 1.9050 ;
      RECT 13.7750 1.5650 13.8650 1.9050 ;
      RECT 14.2950 1.5650 14.3850 1.9050 ;
      RECT 14.8150 1.5650 14.9050 1.9050 ;
      RECT 15.3350 1.5650 15.4250 1.9050 ;
      RECT 15.8550 1.5650 15.9450 1.9050 ;
      RECT 16.3750 1.5650 16.4650 1.9050 ;
      RECT 16.8950 1.5650 16.9850 1.9050 ;
      RECT 17.4150 1.5650 17.5050 1.9050 ;
      RECT 17.9350 1.5650 18.0250 1.9050 ;
      RECT 18.4550 1.5650 18.5450 1.9050 ;
      RECT 18.9750 1.5650 19.0650 1.9050 ;
      RECT 19.4950 1.5650 19.5850 1.9050 ;
      RECT 20.0150 1.5650 20.1050 1.9050 ;
      RECT 20.5350 1.5650 20.6250 1.9050 ;
      RECT 21.0550 1.5650 21.1450 1.9050 ;
      RECT 21.5750 1.5650 21.6650 1.9050 ;
      RECT 22.0950 1.5650 22.1850 1.9050 ;
      RECT 22.6150 1.5650 22.7050 1.9050 ;
      RECT 23.1350 1.5650 23.2250 1.9050 ;
      RECT 23.6550 1.5650 23.7450 1.9050 ;
      RECT 24.1750 1.5650 24.2650 1.9050 ;
      RECT 0.9750 1.2650 24.7850 1.3550 ;
      RECT 24.6950 0.8850 24.7850 1.2650 ;
      RECT 0.7750 0.7950 24.7850 0.8850 ;
      RECT 24.6950 0.4550 24.7850 0.7950 ;
      RECT 0.7750 0.4550 0.8650 0.7950 ;
      RECT 1.2950 0.4550 1.3850 0.7950 ;
      RECT 1.8150 0.4550 1.9050 0.7950 ;
      RECT 2.3350 0.4550 2.4250 0.7950 ;
      RECT 2.8550 0.4550 2.9450 0.7950 ;
      RECT 3.3750 0.4550 3.4650 0.7950 ;
      RECT 3.8950 0.4550 3.9850 0.7950 ;
      RECT 4.4150 0.4550 4.5050 0.7950 ;
      RECT 4.9350 0.4550 5.0250 0.7950 ;
      RECT 5.4550 0.4550 5.5450 0.7950 ;
      RECT 5.9750 0.4550 6.0650 0.7950 ;
      RECT 6.4950 0.4550 6.5850 0.7950 ;
      RECT 7.0150 0.4550 7.1050 0.7950 ;
      RECT 7.5350 0.4550 7.6250 0.7950 ;
      RECT 8.0550 0.4550 8.1450 0.7950 ;
      RECT 8.5750 0.4550 8.6650 0.7950 ;
      RECT 9.0950 0.4550 9.1850 0.7950 ;
      RECT 9.6150 0.4550 9.7050 0.7950 ;
      RECT 10.1350 0.4550 10.2250 0.7950 ;
      RECT 10.6550 0.4550 10.7450 0.7950 ;
      RECT 11.1750 0.4550 11.2650 0.7950 ;
      RECT 11.6950 0.4550 11.7850 0.7950 ;
      RECT 12.2150 0.4550 12.3050 0.7950 ;
      RECT 12.7350 0.4550 12.8250 0.7950 ;
      RECT 13.2550 0.4550 13.3450 0.7950 ;
      RECT 13.7750 0.4550 13.8650 0.7950 ;
      RECT 14.2950 0.4550 14.3850 0.7950 ;
      RECT 14.8150 0.4550 14.9050 0.7950 ;
      RECT 15.3350 0.4550 15.4250 0.7950 ;
      RECT 15.8550 0.4550 15.9450 0.7950 ;
      RECT 16.3750 0.4550 16.4650 0.7950 ;
      RECT 16.8950 0.4550 16.9850 0.7950 ;
      RECT 17.4150 0.4550 17.5050 0.7950 ;
      RECT 17.9350 0.4550 18.0250 0.7950 ;
      RECT 18.4550 0.4550 18.5450 0.7950 ;
      RECT 18.9750 0.4550 19.0650 0.7950 ;
      RECT 19.4950 0.4550 19.5850 0.7950 ;
      RECT 20.0150 0.4550 20.1050 0.7950 ;
      RECT 20.5350 0.4550 20.6250 0.7950 ;
      RECT 21.0550 0.4550 21.1450 0.7950 ;
      RECT 21.5750 0.4550 21.6650 0.7950 ;
      RECT 22.0950 0.4550 22.1850 0.7950 ;
      RECT 22.6150 0.4550 22.7050 0.7950 ;
      RECT 23.1350 0.4550 23.2250 0.7950 ;
      RECT 23.6550 0.4550 23.7450 0.7950 ;
      RECT 24.1750 0.4550 24.2650 0.7950 ;
  END
END FILLCAPTIE128_A12TH

MACRO FILLCAPTIE16_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.5100 1.7700 0.6100 2.0800 ;
        RECT 1.0300 1.7700 1.1300 2.0800 ;
        RECT 1.5500 1.7700 1.6500 2.0800 ;
        RECT 2.0700 1.7700 2.1700 2.0800 ;
        RECT 2.5900 1.7700 2.6900 2.0800 ;
        RECT 0.1350 1.4050 0.2350 2.0800 ;
        RECT 2.9650 1.4050 3.0650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.9750 ;
        RECT 0.5100 0.3200 0.6100 0.6300 ;
        RECT 1.0300 0.3200 1.1300 0.6300 ;
        RECT 1.5500 0.3200 1.6500 0.6300 ;
        RECT 2.0700 0.3200 2.1700 0.6300 ;
        RECT 2.5900 0.3200 2.6900 0.6300 ;
        RECT 2.9650 0.3200 3.0650 0.9750 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.7750 1.4750 2.4250 1.5650 ;
      RECT 2.3350 1.5650 2.4250 1.8850 ;
      RECT 0.7750 1.0050 2.4150 1.0950 ;
      RECT 0.7750 1.5650 0.8650 1.8850 ;
      RECT 0.7750 1.0950 0.8650 1.4750 ;
      RECT 1.2950 1.5650 1.3850 1.9050 ;
      RECT 1.8150 1.5650 1.9050 1.9050 ;
      RECT 0.9750 1.2650 2.6250 1.3550 ;
      RECT 2.5350 0.8850 2.6250 1.2650 ;
      RECT 0.7750 0.7950 2.6250 0.8850 ;
      RECT 0.7750 0.4550 0.8650 0.7950 ;
      RECT 1.2950 0.4550 1.3850 0.7950 ;
      RECT 1.8150 0.4550 1.9050 0.7950 ;
      RECT 2.3350 0.4550 2.4250 0.7950 ;
  END
END FILLCAPTIE16_A12TH

MACRO FILLCAPTIE32_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.5100 1.7700 0.6100 2.0800 ;
        RECT 1.0300 1.7700 1.1300 2.0800 ;
        RECT 1.5500 1.7700 1.6500 2.0800 ;
        RECT 2.0700 1.7700 2.1700 2.0800 ;
        RECT 2.5900 1.7700 2.6900 2.0800 ;
        RECT 3.1100 1.7700 3.2100 2.0800 ;
        RECT 3.6300 1.7700 3.7300 2.0800 ;
        RECT 4.1500 1.7700 4.2500 2.0800 ;
        RECT 4.6700 1.7700 4.7700 2.0800 ;
        RECT 5.1900 1.7700 5.2900 2.0800 ;
        RECT 5.7100 1.7700 5.8100 2.0800 ;
        RECT 0.1350 1.4050 0.2350 2.0800 ;
        RECT 6.1650 1.4050 6.2650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.9750 ;
        RECT 0.5100 0.3200 0.6100 0.6300 ;
        RECT 1.0300 0.3200 1.1300 0.6300 ;
        RECT 1.5500 0.3200 1.6500 0.6300 ;
        RECT 2.0700 0.3200 2.1700 0.6300 ;
        RECT 2.5900 0.3200 2.6900 0.6300 ;
        RECT 3.1100 0.3200 3.2100 0.6300 ;
        RECT 3.6300 0.3200 3.7300 0.6300 ;
        RECT 4.1500 0.3200 4.2500 0.6300 ;
        RECT 4.6700 0.3200 4.7700 0.6300 ;
        RECT 5.1900 0.3200 5.2900 0.6300 ;
        RECT 5.7100 0.3200 5.8100 0.6300 ;
        RECT 6.1650 0.3200 6.2650 0.9750 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.7750 1.4750 5.5450 1.5650 ;
      RECT 5.4550 1.5650 5.5450 1.8850 ;
      RECT 0.7750 1.0050 5.3600 1.0950 ;
      RECT 0.7750 1.5650 0.8650 1.9050 ;
      RECT 0.7750 1.0950 0.8650 1.4750 ;
      RECT 1.2950 1.5650 1.3850 1.9050 ;
      RECT 1.8150 1.5650 1.9050 1.9050 ;
      RECT 2.3350 1.5650 2.4250 1.9050 ;
      RECT 2.8550 1.5650 2.9450 1.9050 ;
      RECT 3.3750 1.5650 3.4650 1.9050 ;
      RECT 3.8950 1.5650 3.9850 1.9050 ;
      RECT 4.4150 1.5650 4.5050 1.9050 ;
      RECT 4.9350 1.5650 5.0250 1.9050 ;
      RECT 0.9750 1.2650 5.6900 1.3550 ;
      RECT 5.6000 0.8850 5.6900 1.2650 ;
      RECT 0.7750 0.7950 5.6900 0.8850 ;
      RECT 5.4550 0.4550 5.5450 0.7950 ;
      RECT 0.7750 0.4550 0.8650 0.7950 ;
      RECT 1.2950 0.4550 1.3850 0.7950 ;
      RECT 1.8150 0.4550 1.9050 0.7950 ;
      RECT 2.3350 0.4550 2.4250 0.7950 ;
      RECT 2.8550 0.4550 2.9450 0.7950 ;
      RECT 3.3750 0.4550 3.4650 0.7950 ;
      RECT 3.8950 0.4550 3.9850 0.7950 ;
      RECT 4.4150 0.4550 4.5050 0.7950 ;
      RECT 4.9350 0.4550 5.0250 0.7950 ;
  END
END FILLCAPTIE32_A12TH

MACRO FILLCAPTIE64_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.8450 2.7200 ;
        RECT 0.5100 1.7700 0.6100 2.0800 ;
        RECT 1.0300 1.7700 1.1300 2.0800 ;
        RECT 1.5500 1.7700 1.6500 2.0800 ;
        RECT 2.0700 1.7700 2.1700 2.0800 ;
        RECT 2.5900 1.7700 2.6900 2.0800 ;
        RECT 3.1100 1.7700 3.2100 2.0800 ;
        RECT 3.6300 1.7700 3.7300 2.0800 ;
        RECT 4.1500 1.7700 4.2500 2.0800 ;
        RECT 4.6700 1.7700 4.7700 2.0800 ;
        RECT 5.1900 1.7700 5.2900 2.0800 ;
        RECT 5.7100 1.7700 5.8100 2.0800 ;
        RECT 6.7500 1.7700 6.8500 2.0800 ;
        RECT 7.2700 1.7700 7.3700 2.0800 ;
        RECT 7.7900 1.7700 7.8900 2.0800 ;
        RECT 8.3100 1.7700 8.4100 2.0800 ;
        RECT 8.8300 1.7700 8.9300 2.0800 ;
        RECT 9.3500 1.7700 9.4500 2.0800 ;
        RECT 9.8700 1.7700 9.9700 2.0800 ;
        RECT 10.3900 1.7700 10.4900 2.0800 ;
        RECT 10.9100 1.7700 11.0100 2.0800 ;
        RECT 11.4300 1.7700 11.5300 2.0800 ;
        RECT 11.9500 1.7700 12.0500 2.0800 ;
        RECT 0.1350 1.4050 0.2350 2.0800 ;
        RECT 12.5650 1.4050 12.6650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.8450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.9750 ;
        RECT 0.5100 0.3200 0.6100 0.6250 ;
        RECT 1.0300 0.3200 1.1300 0.6250 ;
        RECT 1.5500 0.3200 1.6500 0.6250 ;
        RECT 2.0700 0.3200 2.1700 0.6250 ;
        RECT 2.5900 0.3200 2.6900 0.6250 ;
        RECT 3.1100 0.3200 3.2100 0.6250 ;
        RECT 3.6300 0.3200 3.7300 0.6250 ;
        RECT 4.1500 0.3200 4.2500 0.6250 ;
        RECT 4.6700 0.3200 4.7700 0.6250 ;
        RECT 5.1900 0.3200 5.2900 0.6250 ;
        RECT 5.7100 0.3200 5.8100 0.6250 ;
        RECT 6.2300 0.3200 6.3300 0.6250 ;
        RECT 6.7500 0.3200 6.8500 0.6250 ;
        RECT 7.2700 0.3200 7.3700 0.6250 ;
        RECT 7.7900 0.3200 7.8900 0.6250 ;
        RECT 8.3100 0.3200 8.4100 0.6250 ;
        RECT 8.8300 0.3200 8.9300 0.6250 ;
        RECT 9.3500 0.3200 9.4500 0.6250 ;
        RECT 9.8700 0.3200 9.9700 0.6250 ;
        RECT 10.3900 0.3200 10.4900 0.6250 ;
        RECT 10.9100 0.3200 11.0100 0.6250 ;
        RECT 11.4300 0.3200 11.5300 0.6250 ;
        RECT 11.9500 0.3200 12.0500 0.6250 ;
        RECT 12.5650 0.3200 12.6650 0.9750 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.7750 1.4750 12.3050 1.5650 ;
      RECT 12.2150 1.5650 12.3050 1.9050 ;
      RECT 0.7750 1.0050 12.0950 1.0950 ;
      RECT 0.7750 1.5650 0.8650 1.9050 ;
      RECT 0.7750 1.0950 0.8650 1.4750 ;
      RECT 1.2950 1.5650 1.3850 1.9050 ;
      RECT 1.8150 1.5650 1.9050 1.9050 ;
      RECT 2.3350 1.5650 2.4250 1.9050 ;
      RECT 2.8550 1.5650 2.9450 1.9050 ;
      RECT 3.3750 1.5650 3.4650 1.9050 ;
      RECT 3.8950 1.5650 3.9850 1.9050 ;
      RECT 4.4150 1.5650 4.5050 1.9050 ;
      RECT 4.9350 1.5650 5.0250 1.9050 ;
      RECT 5.4550 1.5650 5.5450 1.9050 ;
      RECT 5.9750 1.5650 6.0650 1.9050 ;
      RECT 6.4950 1.5650 6.5850 1.9050 ;
      RECT 7.0150 1.5650 7.1050 1.9050 ;
      RECT 7.5350 1.5650 7.6250 1.9050 ;
      RECT 8.0550 1.5650 8.1450 1.9050 ;
      RECT 8.5750 1.5650 8.6650 1.9050 ;
      RECT 9.0950 1.5650 9.1850 1.9050 ;
      RECT 9.6150 1.5650 9.7050 1.9050 ;
      RECT 10.1350 1.5650 10.2250 1.9050 ;
      RECT 10.6550 1.5650 10.7450 1.9050 ;
      RECT 11.1750 1.5650 11.2650 1.9050 ;
      RECT 11.6950 1.5650 11.7850 1.9050 ;
      RECT 0.9750 1.2650 12.3050 1.3550 ;
      RECT 12.2150 0.8850 12.3050 1.2650 ;
      RECT 0.7750 0.7950 12.3050 0.8850 ;
      RECT 12.2150 0.4350 12.3050 0.7950 ;
      RECT 0.7750 0.4400 0.8650 0.7950 ;
      RECT 1.2950 0.4550 1.3850 0.7950 ;
      RECT 1.8150 0.4550 1.9050 0.7950 ;
      RECT 2.3350 0.4550 2.4250 0.7950 ;
      RECT 2.8550 0.4550 2.9450 0.7950 ;
      RECT 3.3750 0.4550 3.4650 0.7950 ;
      RECT 3.8950 0.4600 3.9850 0.7950 ;
      RECT 4.4150 0.4500 4.5050 0.7950 ;
      RECT 4.9350 0.4550 5.0250 0.7950 ;
      RECT 5.4550 0.4550 5.5450 0.7950 ;
      RECT 5.9750 0.4500 6.0650 0.7950 ;
      RECT 6.4950 0.4550 6.5850 0.7950 ;
      RECT 7.0150 0.4750 7.1050 0.7950 ;
      RECT 7.5350 0.4600 7.6250 0.7950 ;
      RECT 8.0550 0.4550 8.1450 0.7950 ;
      RECT 8.5750 0.4550 8.6650 0.7950 ;
      RECT 9.0950 0.4600 9.1850 0.7950 ;
      RECT 9.6150 0.4600 9.7050 0.7950 ;
      RECT 10.1350 0.4600 10.2250 0.7950 ;
      RECT 10.6550 0.4650 10.7450 0.7950 ;
      RECT 11.1750 0.4650 11.2650 0.7950 ;
      RECT 11.6950 0.4700 11.7850 0.7950 ;
  END
END FILLCAPTIE64_A12TH

MACRO FILLCAPTIE6_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 0.9650 1.3750 1.0650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
        RECT 0.9650 0.3200 1.0650 0.9600 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.3550 1.5100 0.4450 1.8500 ;
      RECT 0.2150 1.4200 0.4450 1.5100 ;
      RECT 0.2150 1.0400 0.3050 1.4200 ;
      RECT 0.0750 0.9500 0.3050 1.0400 ;
      RECT 0.4250 1.2100 0.7050 1.3000 ;
      RECT 0.4250 0.8400 0.5150 1.2100 ;
      RECT 0.3550 0.7500 0.5150 0.8400 ;
      RECT 0.3550 0.4100 0.4450 0.7500 ;
  END
END FILLCAPTIE6_A12TH

MACRO FILLCAPTIE8_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.5100 1.7700 0.6100 2.0800 ;
        RECT 1.0300 1.7700 1.1300 2.0800 ;
        RECT 0.1350 1.3750 0.2350 2.0800 ;
        RECT 1.3650 1.3750 1.4650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.1350 0.3200 0.2350 0.9600 ;
        RECT 0.5100 0.3200 0.6100 0.6300 ;
        RECT 1.0300 0.3200 1.1300 0.6300 ;
        RECT 1.3650 0.3200 1.4650 0.9600 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.7750 1.5100 0.8650 1.8300 ;
      RECT 0.6350 1.4200 0.8650 1.5100 ;
      RECT 0.6350 1.0400 0.7250 1.4200 ;
      RECT 0.4950 0.9500 0.7250 1.0400 ;
      RECT 0.8450 1.2100 1.1150 1.3000 ;
      RECT 0.8450 0.8400 0.9350 1.2100 ;
      RECT 0.7750 0.7500 0.9350 0.8400 ;
      RECT 0.7750 0.4400 0.8650 0.7500 ;
  END
END FILLCAPTIE8_A12TH

MACRO FILLDGCAP128_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 25.6450 2.7200 ;
        RECT 0.9600 0.4700 1.2900 2.0800 ;
        RECT 1.9750 0.4700 2.3050 2.0800 ;
        RECT 2.9900 0.4700 3.3200 2.0800 ;
        RECT 4.0050 0.4700 4.3350 2.0800 ;
        RECT 5.0200 0.4700 5.3500 2.0800 ;
        RECT 6.0350 0.4700 6.3650 2.0800 ;
        RECT 7.0500 0.4700 7.3800 2.0800 ;
        RECT 8.0650 0.4700 8.3950 2.0800 ;
        RECT 9.0800 0.4700 9.4100 2.0800 ;
        RECT 10.0950 0.4700 10.4250 2.0800 ;
        RECT 11.1100 0.4700 11.4400 2.0800 ;
        RECT 12.1250 0.4700 12.4550 2.0800 ;
        RECT 13.1400 0.4700 13.4700 2.0800 ;
        RECT 14.1550 0.4700 14.4850 2.0800 ;
        RECT 15.1700 0.4700 15.5000 2.0800 ;
        RECT 16.1850 0.4700 16.5150 2.0800 ;
        RECT 17.2000 0.4700 17.5300 2.0800 ;
        RECT 18.2150 0.4700 18.5450 2.0800 ;
        RECT 19.2300 0.4700 19.5600 2.0800 ;
        RECT 20.2450 0.4700 20.5750 2.0800 ;
        RECT 21.2600 0.4700 21.5900 2.0800 ;
        RECT 22.2750 0.4700 22.6050 2.0800 ;
        RECT 23.2900 0.4700 23.6200 2.0800 ;
        RECT 24.3050 0.4700 24.6350 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 25.6450 0.3200 ;
        RECT 0.4550 0.3200 0.7850 1.8750 ;
        RECT 1.4700 0.3200 1.8000 1.8750 ;
        RECT 2.4850 0.3200 2.8150 1.8750 ;
        RECT 3.5000 0.3200 3.8300 1.8750 ;
        RECT 4.5150 0.3200 4.8450 1.8750 ;
        RECT 5.5300 0.3200 5.8600 1.8750 ;
        RECT 6.5450 0.3200 6.8750 1.8750 ;
        RECT 7.5600 0.3200 7.8900 1.8750 ;
        RECT 8.5750 0.3200 8.9050 1.8750 ;
        RECT 9.5900 0.3200 9.9200 1.8750 ;
        RECT 10.6050 0.3200 10.9350 1.8750 ;
        RECT 11.6200 0.3200 11.9500 1.8750 ;
        RECT 12.6350 0.3200 12.9650 1.8750 ;
        RECT 13.6500 0.3200 13.9800 1.8750 ;
        RECT 14.6650 0.3200 14.9950 1.8750 ;
        RECT 15.6800 0.3200 16.0100 1.8750 ;
        RECT 16.6950 0.3200 17.0250 1.8750 ;
        RECT 17.7100 0.3200 18.0400 1.8750 ;
        RECT 18.7250 0.3200 19.0550 1.8750 ;
        RECT 19.7400 0.3200 20.0700 1.8750 ;
        RECT 20.7550 0.3200 21.0850 1.8750 ;
        RECT 21.7700 0.3200 22.1000 1.8750 ;
        RECT 22.7850 0.3200 23.1150 1.8750 ;
        RECT 23.8000 0.3200 24.1300 1.8750 ;
        RECT 24.8150 0.3200 25.1450 1.8750 ;
    END
  END VSS
END FILLDGCAP128_A12TH

MACRO FILLDGCAP12_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.9900 0.4800 1.4100 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.4900 0.3200 0.7500 1.8750 ;
        RECT 1.6500 0.3200 1.9100 1.8750 ;
    END
  END VSS
END FILLDGCAP12_A12TH

MACRO FILLDGCAP16_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.9250 0.5000 1.2950 2.0800 ;
        RECT 1.9050 0.5000 2.2750 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.4550 0.3200 0.7850 1.8750 ;
        RECT 1.4350 0.3200 1.7650 1.8600 ;
        RECT 2.4150 0.3200 2.7450 1.8750 ;
    END
  END VSS
END FILLDGCAP16_A12TH

MACRO FILLDGCAP32_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.9750 0.4700 1.3050 2.0800 ;
        RECT 2.0050 0.4700 2.3350 2.0800 ;
        RECT 3.0350 0.4700 3.3650 2.0800 ;
        RECT 4.0650 0.4700 4.3950 2.0800 ;
        RECT 5.0950 0.4700 5.4250 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.4550 0.3200 0.7900 1.7600 ;
        RECT 1.4900 0.3200 1.8200 1.8750 ;
        RECT 2.5200 0.3200 2.8500 1.8750 ;
        RECT 3.5500 0.3200 3.8800 1.8750 ;
        RECT 4.5800 0.3200 4.9100 1.8750 ;
        RECT 5.6100 0.3200 5.9400 1.8750 ;
        RECT 0.4600 1.7600 0.7900 1.8750 ;
    END
  END VSS
END FILLDGCAP32_A12TH

MACRO FILLDGCAP64_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.8450 2.7200 ;
        RECT 0.9850 0.4700 1.3150 2.0800 ;
        RECT 2.0350 0.4700 2.3650 2.0800 ;
        RECT 3.0850 0.4700 3.4150 2.0800 ;
        RECT 4.1350 0.4700 4.4650 2.0800 ;
        RECT 5.1850 0.4700 5.5150 2.0800 ;
        RECT 6.2350 0.4700 6.5650 2.0800 ;
        RECT 7.2850 0.4700 7.6150 2.0800 ;
        RECT 8.3350 0.4700 8.6650 2.0800 ;
        RECT 9.3850 0.4700 9.7150 2.0800 ;
        RECT 10.4350 0.4700 10.7650 2.0800 ;
        RECT 11.4850 0.4700 11.8150 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.8450 0.3200 ;
        RECT 0.4600 0.3200 0.7900 1.8750 ;
        RECT 1.5100 0.3200 1.8400 1.8750 ;
        RECT 2.5600 0.3200 2.8900 1.8750 ;
        RECT 3.6100 0.3200 3.9400 1.8750 ;
        RECT 4.6600 0.3200 4.9900 1.8750 ;
        RECT 5.7100 0.3200 6.0400 1.8750 ;
        RECT 6.7600 0.3200 7.0900 1.8750 ;
        RECT 7.8100 0.3200 8.1400 1.8750 ;
        RECT 8.8600 0.3200 9.1900 1.8750 ;
        RECT 9.9100 0.3200 10.2400 1.8750 ;
        RECT 10.9600 0.3200 11.2900 1.8750 ;
        RECT 12.0100 0.3200 12.3400 1.8750 ;
    END
  END VSS
END FILLDGCAP64_A12TH

MACRO FILLDGCAPTIE128_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 25.6450 2.7200 ;
        RECT 0.1250 1.4250 0.2550 2.0800 ;
        RECT 25.3450 1.4250 25.4750 2.0800 ;
        RECT 1.1950 0.4700 1.5250 2.0800 ;
        RECT 2.2350 0.4700 2.5650 2.0800 ;
        RECT 3.2750 0.4700 3.6050 2.0800 ;
        RECT 4.3150 0.4700 4.6450 2.0800 ;
        RECT 5.3550 0.4700 5.6850 2.0800 ;
        RECT 6.3950 0.4700 6.7250 2.0800 ;
        RECT 7.4350 0.4700 7.7650 2.0800 ;
        RECT 8.4750 0.4700 8.8050 2.0800 ;
        RECT 9.5150 0.4700 9.8450 2.0800 ;
        RECT 10.5550 0.4700 10.8850 2.0800 ;
        RECT 11.5950 0.4700 11.9250 2.0800 ;
        RECT 12.6350 0.4700 12.9650 2.0800 ;
        RECT 13.6750 0.4700 14.0050 2.0800 ;
        RECT 14.7150 0.4700 15.0450 2.0800 ;
        RECT 15.7550 0.4700 16.0850 2.0800 ;
        RECT 16.7950 0.4700 17.1250 2.0800 ;
        RECT 17.8350 0.4700 18.1650 2.0800 ;
        RECT 18.8750 0.4700 19.2050 2.0800 ;
        RECT 19.9150 0.4700 20.2450 2.0800 ;
        RECT 20.9550 0.4700 21.2850 2.0800 ;
        RECT 21.9950 0.4700 22.3250 2.0800 ;
        RECT 23.0350 0.4700 23.3650 2.0800 ;
        RECT 24.0750 0.4700 24.4050 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 25.6450 0.3200 ;
        RECT 0.1250 0.3200 0.2550 0.9000 ;
        RECT 0.7550 0.3200 0.9250 1.8750 ;
        RECT 1.7950 0.3200 1.9650 1.8750 ;
        RECT 2.8350 0.3200 3.0050 1.8750 ;
        RECT 3.8750 0.3200 4.0450 1.8750 ;
        RECT 4.9150 0.3200 5.0850 1.8750 ;
        RECT 5.9550 0.3200 6.1250 1.8750 ;
        RECT 6.9950 0.3200 7.1650 1.8750 ;
        RECT 8.0350 0.3200 8.2050 1.8750 ;
        RECT 9.0750 0.3200 9.2450 1.8750 ;
        RECT 10.1150 0.3200 10.2850 1.8750 ;
        RECT 11.1550 0.3200 11.3250 1.8750 ;
        RECT 12.1950 0.3200 12.3650 1.8750 ;
        RECT 13.2350 0.3200 13.4050 1.8750 ;
        RECT 14.2750 0.3200 14.4450 1.8750 ;
        RECT 15.3150 0.3200 15.4850 1.8750 ;
        RECT 16.3550 0.3200 16.5250 1.8750 ;
        RECT 17.3950 0.3200 17.5650 1.8750 ;
        RECT 18.4350 0.3200 18.6050 1.8750 ;
        RECT 19.4750 0.3200 19.6450 1.8750 ;
        RECT 20.5150 0.3200 20.6850 1.8750 ;
        RECT 21.5550 0.3200 21.7250 1.8750 ;
        RECT 22.5950 0.3200 22.7650 1.8750 ;
        RECT 23.6350 0.3200 23.8050 1.8750 ;
        RECT 24.6750 0.3200 24.8450 1.8750 ;
        RECT 25.3450 0.3200 25.4750 0.9000 ;
    END
  END VSS
END FILLDGCAPTIE128_A12TH

MACRO FILLDGCAPTIE12_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.1250 1.4250 0.2550 2.0800 ;
        RECT 2.1450 1.4250 2.2750 2.0800 ;
        RECT 1.0350 0.4700 1.3650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1250 0.3200 0.2550 0.9000 ;
        RECT 0.7450 0.3200 0.8750 1.8750 ;
        RECT 1.5250 0.3200 1.6550 1.8750 ;
        RECT 2.1450 0.3200 2.2750 0.9000 ;
    END
  END VSS
END FILLDGCAPTIE12_A12TH

MACRO FILLDGCAPTIE16_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.1250 1.4250 0.2550 2.0800 ;
        RECT 2.9450 1.4250 3.0750 2.0800 ;
        RECT 1.1150 0.4700 1.4450 2.0800 ;
        RECT 1.7550 0.4700 2.0850 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.1250 0.3200 0.2550 0.9000 ;
        RECT 0.7450 0.3200 0.8750 1.8750 ;
        RECT 2.3250 0.3200 2.4550 1.8750 ;
        RECT 2.9450 0.3200 3.0750 0.9000 ;
    END
  END VSS
END FILLDGCAPTIE16_A12TH

MACRO FILLDGCAPTIE32_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.1250 1.4250 0.2550 2.0800 ;
        RECT 6.1450 1.4250 6.2750 2.0800 ;
        RECT 1.2250 0.4700 1.5950 2.0800 ;
        RECT 2.4200 0.4700 2.7900 2.0800 ;
        RECT 3.6150 0.4700 3.9850 2.0800 ;
        RECT 4.8100 0.4700 5.1800 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.1250 0.3200 0.2550 0.9000 ;
        RECT 0.7250 0.3200 0.8950 1.8650 ;
        RECT 1.9200 0.3200 2.0900 1.8650 ;
        RECT 3.1150 0.3200 3.2850 1.8650 ;
        RECT 4.3100 0.3200 4.4800 1.8650 ;
        RECT 5.5050 0.3200 5.6750 1.8650 ;
        RECT 6.1450 0.3200 6.2750 0.9000 ;
    END
  END VSS
END FILLDGCAPTIE32_A12TH

MACRO FILLDGCAPTIE64_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.8450 2.7200 ;
        RECT 0.1250 1.4250 0.2550 2.0800 ;
        RECT 12.5450 1.4250 12.6750 2.0800 ;
        RECT 1.1400 0.4700 1.5100 2.0800 ;
        RECT 2.1550 0.4700 2.5250 2.0800 ;
        RECT 3.1700 0.4700 3.5400 2.0800 ;
        RECT 4.1850 0.4700 4.5550 2.0800 ;
        RECT 5.2000 0.4700 5.5700 2.0800 ;
        RECT 6.2150 0.4700 6.5850 2.0800 ;
        RECT 7.2300 0.4700 7.6000 2.0800 ;
        RECT 8.2450 0.4700 8.6150 2.0800 ;
        RECT 9.2600 0.4700 9.6300 2.0800 ;
        RECT 10.2750 0.4700 10.6450 2.0800 ;
        RECT 11.2900 0.4700 11.6600 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.8450 0.3200 ;
        RECT 0.1250 0.3200 0.2550 0.9000 ;
        RECT 0.7300 0.3200 0.9000 1.8750 ;
        RECT 1.7450 0.3200 1.9150 1.8750 ;
        RECT 2.7600 0.3200 2.9300 1.8750 ;
        RECT 3.7750 0.3200 3.9450 1.8750 ;
        RECT 4.7900 0.3200 4.9600 1.8750 ;
        RECT 5.8050 0.3200 5.9750 1.8750 ;
        RECT 6.8200 0.3200 6.9900 1.8750 ;
        RECT 7.8350 0.3200 8.0050 1.8750 ;
        RECT 8.8500 0.3200 9.0200 1.8750 ;
        RECT 9.8650 0.3200 10.0350 1.8750 ;
        RECT 10.8800 0.3200 11.0500 1.8750 ;
        RECT 11.8950 0.3200 12.0650 1.8750 ;
        RECT 12.5450 0.3200 12.6750 0.9000 ;
    END
  END VSS
END FILLDGCAPTIE64_A12TH

MACRO FILLTIE128_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 25.6450 2.7200 ;
        RECT 19.3200 1.9900 19.4900 2.0800 ;
        RECT 19.7200 1.9900 19.8900 2.0800 ;
        RECT 20.1200 1.9900 20.2900 2.0800 ;
        RECT 20.5150 1.9900 20.6850 2.0800 ;
        RECT 20.9200 1.9900 21.0900 2.0800 ;
        RECT 21.3200 1.9900 21.4900 2.0800 ;
        RECT 21.7200 1.9900 21.8900 2.0800 ;
        RECT 22.1200 1.9900 22.2900 2.0800 ;
        RECT 22.5200 1.9900 22.6900 2.0800 ;
        RECT 22.9200 1.9900 23.0900 2.0800 ;
        RECT 23.3200 1.9900 23.4900 2.0800 ;
        RECT 23.7200 1.9900 23.8900 2.0800 ;
        RECT 24.1200 1.9900 24.2900 2.0800 ;
        RECT 24.5200 1.9900 24.6900 2.0800 ;
        RECT 24.9200 1.9900 25.0900 2.0800 ;
        RECT 25.3500 1.5050 25.4500 2.0800 ;
        RECT 12.9200 1.9900 13.0900 2.0800 ;
        RECT 13.3200 1.9900 13.4900 2.0800 ;
        RECT 13.7200 1.9900 13.8900 2.0800 ;
        RECT 14.1200 1.9900 14.2900 2.0800 ;
        RECT 14.5200 1.9900 14.6900 2.0800 ;
        RECT 14.9150 1.9900 15.0850 2.0800 ;
        RECT 15.3200 1.9900 15.4900 2.0800 ;
        RECT 15.7200 1.9900 15.8900 2.0800 ;
        RECT 16.1200 1.9900 16.2900 2.0800 ;
        RECT 16.5200 1.9900 16.6900 2.0800 ;
        RECT 16.9200 1.9900 17.0900 2.0800 ;
        RECT 17.3200 1.9900 17.4900 2.0800 ;
        RECT 17.7200 1.9900 17.8900 2.0800 ;
        RECT 18.1150 1.9900 18.2850 2.0800 ;
        RECT 18.5200 1.9900 18.6900 2.0800 ;
        RECT 18.9200 1.9900 19.0900 2.0800 ;
        RECT 6.5200 1.9900 6.6900 2.0800 ;
        RECT 6.9200 1.9900 7.0900 2.0800 ;
        RECT 7.3200 1.9900 7.4900 2.0800 ;
        RECT 7.7200 1.9900 7.8900 2.0800 ;
        RECT 8.1200 1.9900 8.2900 2.0800 ;
        RECT 8.5150 1.9900 8.6850 2.0800 ;
        RECT 8.9200 1.9900 9.0900 2.0800 ;
        RECT 9.3200 1.9900 9.4900 2.0800 ;
        RECT 9.7200 1.9900 9.8900 2.0800 ;
        RECT 10.1200 1.9900 10.2900 2.0800 ;
        RECT 10.5200 1.9900 10.6900 2.0800 ;
        RECT 10.9200 1.9900 11.0900 2.0800 ;
        RECT 11.3200 1.9900 11.4900 2.0800 ;
        RECT 11.7200 1.9900 11.8900 2.0800 ;
        RECT 12.1200 1.9900 12.2900 2.0800 ;
        RECT 12.5150 1.9900 12.6850 2.0800 ;
        RECT 0.5150 1.9900 0.6850 2.0800 ;
        RECT 0.9200 1.9900 1.0900 2.0800 ;
        RECT 1.3200 1.9900 1.4900 2.0800 ;
        RECT 1.7200 1.9900 1.8900 2.0800 ;
        RECT 2.1200 1.9900 2.2900 2.0800 ;
        RECT 2.5200 1.9900 2.6900 2.0800 ;
        RECT 2.9150 1.9900 3.0850 2.0800 ;
        RECT 3.3200 1.9900 3.4900 2.0800 ;
        RECT 3.7200 1.9900 3.8900 2.0800 ;
        RECT 4.1200 1.9900 4.2900 2.0800 ;
        RECT 4.5200 1.9900 4.6900 2.0800 ;
        RECT 4.9200 1.9900 5.0900 2.0800 ;
        RECT 5.3200 1.9900 5.4900 2.0800 ;
        RECT 5.7200 1.9900 5.8900 2.0800 ;
        RECT 6.1150 1.9900 6.2850 2.0800 ;
        RECT 0.1500 1.5050 0.2500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 25.6450 0.3200 ;
        RECT 25.3500 0.3200 25.4500 0.8550 ;
        RECT 19.3150 0.3200 19.4850 0.4100 ;
        RECT 19.7150 0.3200 19.8850 0.4100 ;
        RECT 20.1150 0.3200 20.2850 0.4100 ;
        RECT 20.5150 0.3200 20.6850 0.4100 ;
        RECT 20.9150 0.3200 21.0850 0.4100 ;
        RECT 21.3150 0.3200 21.4850 0.4100 ;
        RECT 21.7150 0.3200 21.8850 0.4100 ;
        RECT 22.1150 0.3200 22.2850 0.4100 ;
        RECT 22.5150 0.3200 22.6850 0.4100 ;
        RECT 22.9150 0.3200 23.0850 0.4100 ;
        RECT 23.3150 0.3200 23.4850 0.4100 ;
        RECT 23.7150 0.3200 23.8850 0.4100 ;
        RECT 24.1150 0.3200 24.2850 0.4100 ;
        RECT 24.5150 0.3200 24.6850 0.4100 ;
        RECT 24.9150 0.3200 25.0850 0.4100 ;
        RECT 12.9150 0.3200 13.0850 0.4100 ;
        RECT 13.3150 0.3200 13.4850 0.4100 ;
        RECT 13.7150 0.3200 13.8850 0.4100 ;
        RECT 14.1150 0.3200 14.2850 0.4100 ;
        RECT 14.5150 0.3200 14.6850 0.4100 ;
        RECT 14.9150 0.3200 15.0850 0.4100 ;
        RECT 15.3150 0.3200 15.4850 0.4100 ;
        RECT 15.7150 0.3200 15.8850 0.4100 ;
        RECT 16.1150 0.3200 16.2850 0.4100 ;
        RECT 16.5150 0.3200 16.6850 0.4100 ;
        RECT 16.9150 0.3200 17.0850 0.4100 ;
        RECT 17.3150 0.3200 17.4850 0.4100 ;
        RECT 17.7150 0.3200 17.8850 0.4100 ;
        RECT 18.1150 0.3200 18.2850 0.4100 ;
        RECT 18.5150 0.3200 18.6850 0.4100 ;
        RECT 18.9150 0.3200 19.0850 0.4100 ;
        RECT 6.5150 0.3200 6.6850 0.4100 ;
        RECT 6.9150 0.3200 7.0850 0.4100 ;
        RECT 7.3150 0.3200 7.4850 0.4100 ;
        RECT 7.7150 0.3200 7.8850 0.4100 ;
        RECT 8.1150 0.3200 8.2850 0.4100 ;
        RECT 8.5150 0.3200 8.6850 0.4100 ;
        RECT 8.9150 0.3200 9.0850 0.4100 ;
        RECT 9.3150 0.3200 9.4850 0.4100 ;
        RECT 9.7150 0.3200 9.8850 0.4100 ;
        RECT 10.1150 0.3200 10.2850 0.4100 ;
        RECT 10.5150 0.3200 10.6850 0.4100 ;
        RECT 10.9150 0.3200 11.0850 0.4100 ;
        RECT 11.3150 0.3200 11.4850 0.4100 ;
        RECT 11.7150 0.3200 11.8850 0.4100 ;
        RECT 12.1150 0.3200 12.2850 0.4100 ;
        RECT 12.5150 0.3200 12.6850 0.4100 ;
        RECT 0.1500 0.3200 0.2500 0.8550 ;
        RECT 0.5150 0.3200 0.6850 0.4100 ;
        RECT 0.9150 0.3200 1.0850 0.4100 ;
        RECT 1.3150 0.3200 1.4850 0.4100 ;
        RECT 1.7150 0.3200 1.8850 0.4100 ;
        RECT 2.1150 0.3200 2.2850 0.4100 ;
        RECT 2.5150 0.3200 2.6850 0.4100 ;
        RECT 2.9150 0.3200 3.0850 0.4100 ;
        RECT 3.3150 0.3200 3.4850 0.4100 ;
        RECT 3.7150 0.3200 3.8850 0.4100 ;
        RECT 4.1150 0.3200 4.2850 0.4100 ;
        RECT 4.5150 0.3200 4.6850 0.4100 ;
        RECT 4.9150 0.3200 5.0850 0.4100 ;
        RECT 5.3150 0.3200 5.4850 0.4100 ;
        RECT 5.7150 0.3200 5.8850 0.4100 ;
        RECT 6.1150 0.3200 6.2850 0.4100 ;
    END
  END VSS
END FILLTIE128_A12TH

MACRO DLY4_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.5350 1.7700 0.6350 2.0800 ;
        RECT 1.7050 1.7700 1.8050 2.0800 ;
        RECT 1.9650 1.7700 2.0650 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.5350 0.3200 0.6350 0.6350 ;
        RECT 1.7050 0.3200 1.8050 0.6350 ;
        RECT 1.9650 0.3200 2.0650 0.6350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9300 2.3500 1.5450 ;
        RECT 2.2250 1.5450 2.3500 1.6450 ;
        RECT 2.2250 0.8100 2.3500 0.9300 ;
        RECT 2.2250 1.6450 2.3250 1.9750 ;
        RECT 2.2250 0.4900 2.3250 0.8100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1250 1.0500 0.5500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5450 0.8850 1.6450 ;
      RECT 0.7850 0.9000 0.8850 1.5450 ;
      RECT 0.0750 0.8000 0.8850 0.9000 ;
      RECT 0.0750 1.6450 0.1750 1.9750 ;
      RECT 0.0750 0.5350 0.1750 0.8000 ;
      RECT 0.9950 1.1500 1.0950 1.9900 ;
      RECT 0.9950 1.0500 1.6550 1.1500 ;
      RECT 0.9950 0.5350 1.0950 1.0500 ;
      RECT 1.8550 1.0550 2.0800 1.1550 ;
      RECT 1.2450 1.5500 1.3450 1.9900 ;
      RECT 1.2450 0.5350 1.3450 0.8450 ;
      RECT 1.2450 1.4500 1.9550 1.5500 ;
      RECT 1.8550 1.1550 1.9550 1.4500 ;
      RECT 1.8550 0.9450 1.9550 1.0550 ;
      RECT 1.2450 0.8450 1.9550 0.9450 ;
  END
END DLY4_X1M_A12TH

MACRO DLY4_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.5750 1.7700 0.6750 2.0800 ;
        RECT 1.8250 1.7700 1.9250 2.0800 ;
        RECT 2.0850 1.7700 2.1850 2.0800 ;
        RECT 2.6050 1.7700 2.7050 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.5750 0.3200 0.6750 0.6350 ;
        RECT 1.8250 0.3200 1.9250 0.6350 ;
        RECT 2.0850 0.3200 2.1850 0.6350 ;
        RECT 2.6050 0.3200 2.7050 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1500 1.0500 0.5900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1584 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9300 2.5500 1.5450 ;
        RECT 2.3450 1.5450 2.5500 1.6450 ;
        RECT 2.3450 0.8100 2.5500 0.9300 ;
        RECT 2.3450 1.6450 2.4450 1.9750 ;
        RECT 2.3450 0.4900 2.4450 0.8100 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5450 0.9250 1.6450 ;
      RECT 0.8250 0.9000 0.9250 1.5450 ;
      RECT 0.0750 0.8000 0.9250 0.9000 ;
      RECT 0.0750 1.6450 0.1750 1.9750 ;
      RECT 0.0750 0.5350 0.1750 0.8000 ;
      RECT 1.0750 1.1500 1.1750 1.8900 ;
      RECT 1.0750 1.0500 1.7750 1.1500 ;
      RECT 1.0750 0.5350 1.1750 1.0500 ;
      RECT 1.9750 1.0550 2.3600 1.1550 ;
      RECT 1.3250 1.5500 1.4250 1.8900 ;
      RECT 1.3250 0.5350 1.4250 0.8450 ;
      RECT 1.3250 1.4500 2.0750 1.5500 ;
      RECT 1.9750 1.1550 2.0750 1.4500 ;
      RECT 1.9750 0.9450 2.0750 1.0550 ;
      RECT 1.3250 0.8450 2.0750 0.9450 ;
  END
END DLY4_X2M_A12TH

MACRO DLY4_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0750 1.7700 0.1750 2.0800 ;
        RECT 1.0450 1.7700 1.1450 2.0800 ;
        RECT 2.0250 1.7700 2.1250 2.0800 ;
        RECT 2.2750 1.7700 2.3750 2.0800 ;
        RECT 3.2550 1.7700 3.3550 2.0800 ;
        RECT 3.5150 1.7700 3.6150 2.0800 ;
        RECT 3.7750 1.7700 3.8750 2.0800 ;
        RECT 4.2950 1.7700 4.3950 2.0800 ;
        RECT 4.8150 1.7700 4.9150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.9500 4.7500 1.2500 ;
        RECT 4.0350 1.2500 4.7500 1.3500 ;
        RECT 4.0350 0.8500 4.7500 0.9500 ;
        RECT 4.0350 1.3500 4.1350 1.7200 ;
        RECT 4.5550 1.3500 4.6550 1.7200 ;
        RECT 4.0350 0.4900 4.1350 0.8500 ;
        RECT 4.5550 0.4900 4.6550 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0500 0.9650 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6350 ;
        RECT 1.0450 0.3200 1.1450 0.6350 ;
        RECT 2.0250 0.3200 2.1250 0.6350 ;
        RECT 2.2750 0.3200 2.3750 0.6350 ;
        RECT 3.2550 0.3200 3.3550 0.6350 ;
        RECT 3.5150 0.3200 3.6150 0.6350 ;
        RECT 3.7750 0.3200 3.8750 0.6350 ;
        RECT 4.2950 0.3200 4.3950 0.6350 ;
        RECT 4.8150 0.3200 4.9150 0.6350 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.5550 1.4500 1.3950 1.5500 ;
      RECT 1.2950 1.1550 1.3950 1.4500 ;
      RECT 1.2950 1.0550 1.8800 1.1550 ;
      RECT 1.2950 0.9000 1.3950 1.0550 ;
      RECT 0.5550 0.8000 1.3950 0.9000 ;
      RECT 0.5550 1.5500 0.6550 1.9200 ;
      RECT 0.5550 0.4300 0.6550 0.8000 ;
      RECT 2.0100 1.0500 3.2150 1.1500 ;
      RECT 1.5350 1.5500 1.6350 1.8900 ;
      RECT 1.5350 0.4300 1.6350 0.7400 ;
      RECT 1.5350 1.4500 2.1100 1.5500 ;
      RECT 2.0100 1.1500 2.1100 1.4500 ;
      RECT 2.0100 0.8400 2.1100 1.0500 ;
      RECT 1.5350 0.7400 2.1100 0.8400 ;
      RECT 3.4050 1.0550 4.5050 1.1550 ;
      RECT 2.7650 1.5500 2.8650 1.8900 ;
      RECT 2.7650 0.4300 2.8650 0.8450 ;
      RECT 2.7650 1.4500 3.5050 1.5500 ;
      RECT 3.4050 1.1550 3.5050 1.4500 ;
      RECT 3.4050 0.9450 3.5050 1.0550 ;
      RECT 2.7650 0.8450 3.5050 0.9450 ;
  END
END DLY4_X4M_A12TH

MACRO EDFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.4000 0.3200 0.5200 0.7600 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9150 0.7500 1.3400 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8600 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 1.1550 6.2500 1.3900 ;
        RECT 6.1200 0.9650 6.2500 1.1550 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2250 1.4050 5.4800 1.6850 ;
        RECT 5.3900 0.7850 5.4800 1.4050 ;
    END
    ANTENNADIFFAREA 0.1233 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.3550 1.9950 0.5650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6900 1.5250 0.9300 1.6150 ;
      RECT 0.8400 0.7450 0.9300 1.5250 ;
      RECT 0.6750 0.6550 0.9300 0.7450 ;
      RECT 0.3050 1.7650 1.0600 1.8550 ;
      RECT 0.3050 1.7050 0.3950 1.7650 ;
      RECT 0.0550 1.6150 0.3950 1.7050 ;
      RECT 0.0550 0.7150 0.1450 1.6150 ;
      RECT 0.0550 0.6250 0.2450 0.7150 ;
      RECT 1.0200 0.5700 1.1100 1.6500 ;
      RECT 1.0200 0.4800 1.7350 0.5700 ;
      RECT 1.6450 0.5700 1.7350 1.3350 ;
      RECT 1.8450 0.6050 1.9450 1.6350 ;
      RECT 2.0800 1.4700 2.3050 1.5600 ;
      RECT 2.2150 0.7700 2.3050 1.4700 ;
      RECT 2.2150 0.6800 3.0150 0.7700 ;
      RECT 2.9250 0.7700 3.0150 1.3150 ;
      RECT 2.5800 1.4700 3.2800 1.5600 ;
      RECT 2.5800 1.0500 2.6700 1.4700 ;
      RECT 3.1900 0.7700 3.2800 1.4700 ;
      RECT 3.1100 0.6800 3.2800 0.7700 ;
      RECT 3.3900 1.4700 3.9250 1.5600 ;
      RECT 3.8350 0.7700 3.9250 1.4700 ;
      RECT 3.5500 0.6800 4.3050 0.7700 ;
      RECT 4.2150 0.7700 4.3050 0.9500 ;
      RECT 4.2150 0.9500 4.3800 1.1650 ;
      RECT 1.3200 1.8300 2.1250 1.9200 ;
      RECT 2.0350 1.7400 2.1250 1.8300 ;
      RECT 1.3200 0.7500 1.4100 1.8300 ;
      RECT 2.0350 1.6500 4.8700 1.7400 ;
      RECT 1.2200 0.6600 1.4100 0.7500 ;
      RECT 4.7800 0.9500 4.8700 1.6500 ;
      RECT 4.6850 0.8600 4.8700 0.9500 ;
      RECT 4.3950 0.6800 5.2750 0.7700 ;
      RECT 5.1850 0.7700 5.2750 1.2700 ;
      RECT 4.0150 1.4200 4.5750 1.5100 ;
      RECT 4.4850 1.2500 4.5750 1.4200 ;
      RECT 4.0150 1.0250 4.1050 1.4200 ;
      RECT 4.4850 1.0400 4.6450 1.2500 ;
      RECT 4.4850 0.7700 4.5750 1.0400 ;
      RECT 2.0350 0.4800 5.7100 0.5700 ;
      RECT 5.5800 0.5700 5.7100 0.6750 ;
      RECT 5.6200 0.6750 5.7100 1.7200 ;
      RECT 3.3700 1.2700 3.7350 1.3600 ;
      RECT 3.3700 0.5700 3.4600 1.2700 ;
      RECT 2.0350 0.5700 2.1250 1.3600 ;
      RECT 2.3550 0.4100 2.5250 0.4800 ;
      RECT 5.8000 1.6600 6.3200 1.7500 ;
      RECT 6.2300 1.5700 6.3200 1.6600 ;
      RECT 5.8000 0.5650 6.3200 0.6550 ;
      RECT 6.2300 0.4850 6.3200 0.5650 ;
      RECT 2.2750 1.8300 5.8900 1.9200 ;
      RECT 5.8000 1.7500 5.8900 1.8300 ;
      RECT 5.8000 0.6550 5.8900 1.6600 ;
  END
END EDFFQN_X0P5M_A12TH

MACRO EDFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.4000 0.3200 0.5200 0.7150 ;
        RECT 4.9650 0.3200 5.1350 0.3550 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8250 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8350 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0200 0.9650 6.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2450 1.4050 5.4150 1.6850 ;
        RECT 5.3150 0.6900 5.4150 1.4050 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 0.4100 1.9250 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6900 1.4500 0.9500 1.5400 ;
      RECT 0.8500 0.6650 0.9500 1.4500 ;
      RECT 0.6750 0.5750 0.9500 0.6650 ;
      RECT 0.3050 1.7400 1.0600 1.8300 ;
      RECT 0.3050 1.6150 0.3950 1.7400 ;
      RECT 0.0550 1.5250 0.3950 1.6150 ;
      RECT 0.0550 0.6650 0.1450 1.5250 ;
      RECT 0.0550 0.5750 0.2450 0.6650 ;
      RECT 1.0400 0.5700 1.1300 1.5700 ;
      RECT 1.0400 0.4800 1.7750 0.5700 ;
      RECT 1.6850 0.5700 1.7750 1.3350 ;
      RECT 1.8850 0.5250 1.9850 1.6600 ;
      RECT 2.1200 1.4700 2.3450 1.5600 ;
      RECT 2.2550 0.7700 2.3450 1.4700 ;
      RECT 2.2550 0.6800 3.0200 0.7700 ;
      RECT 2.9300 0.7700 3.0200 1.3250 ;
      RECT 2.6200 1.4700 3.2800 1.5600 ;
      RECT 2.6200 1.0600 2.7100 1.4700 ;
      RECT 3.1900 0.7700 3.2800 1.4700 ;
      RECT 3.1100 0.6800 3.2800 0.7700 ;
      RECT 3.3900 1.4700 3.9250 1.5600 ;
      RECT 3.8350 0.7700 3.9250 1.4700 ;
      RECT 3.5500 0.6800 4.3050 0.7700 ;
      RECT 4.2150 0.7700 4.3050 0.9550 ;
      RECT 4.2150 0.9550 4.3800 1.1650 ;
      RECT 1.3400 1.7700 2.1650 1.8600 ;
      RECT 2.0750 1.7400 2.1650 1.7700 ;
      RECT 1.3400 0.7500 1.4300 1.7700 ;
      RECT 2.0750 1.6500 4.8800 1.7400 ;
      RECT 1.2400 0.6600 1.4300 0.7500 ;
      RECT 4.7900 0.9500 4.8800 1.6500 ;
      RECT 4.6950 0.8600 4.8800 0.9500 ;
      RECT 4.0150 1.4200 4.5750 1.5100 ;
      RECT 4.4850 1.2100 4.5750 1.4200 ;
      RECT 4.0150 1.0250 4.1050 1.4200 ;
      RECT 4.4850 1.0400 4.6800 1.2100 ;
      RECT 4.4850 0.7700 4.5750 1.0400 ;
      RECT 4.3950 0.6800 5.2200 0.7700 ;
      RECT 5.1300 0.7700 5.2200 1.2200 ;
      RECT 2.0750 0.4800 5.6600 0.5700 ;
      RECT 5.5700 0.5700 5.6600 1.7200 ;
      RECT 3.3700 1.2700 3.7350 1.3600 ;
      RECT 3.3700 0.5700 3.4600 1.2700 ;
      RECT 2.0750 0.5700 2.1650 1.3600 ;
      RECT 2.3950 0.4100 2.5650 0.4800 ;
      RECT 5.7650 1.6500 6.3400 1.7400 ;
      RECT 5.7650 0.5550 6.3400 0.6450 ;
      RECT 2.2950 1.8300 5.8550 1.9200 ;
      RECT 5.7650 1.7400 5.8550 1.8300 ;
      RECT 5.7650 0.6450 5.8550 1.6500 ;
  END
END EDFFQN_X1M_A12TH

MACRO EDFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.4000 0.3200 0.5200 0.6950 ;
        RECT 3.8800 0.3200 4.2500 0.3600 ;
        RECT 4.9450 0.3200 5.1150 0.3550 ;
        RECT 5.5050 0.3200 5.6750 0.3550 ;
        RECT 6.0800 0.3200 6.2500 0.5000 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2850 1.2500 5.6000 1.3500 ;
        RECT 5.2850 1.3500 5.3750 1.7200 ;
        RECT 5.5000 0.8450 5.6000 1.2500 ;
        RECT 5.2300 0.7450 5.6000 0.8450 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2500 0.9650 6.4100 1.3900 ;
    END
    ANTENNAGATEAREA 0.033 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 0.8450 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0528 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8350 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END E

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 4.1100 2.0200 4.2800 2.0800 ;
        RECT 0.4100 1.9250 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6900 1.4500 0.9500 1.5400 ;
      RECT 0.8500 0.6650 0.9500 1.4500 ;
      RECT 0.6750 0.5750 0.9500 0.6650 ;
      RECT 0.0500 1.7400 1.0600 1.8300 ;
      RECT 0.0500 0.6650 0.1400 1.7400 ;
      RECT 0.0500 0.5750 0.2450 0.6650 ;
      RECT 1.0400 0.5700 1.1300 1.5700 ;
      RECT 1.0400 0.4800 1.7750 0.5700 ;
      RECT 1.6850 0.5700 1.7750 1.3150 ;
      RECT 1.8850 0.5250 1.9850 1.6600 ;
      RECT 2.1200 1.4700 2.3450 1.5600 ;
      RECT 2.2550 0.7700 2.3450 1.4700 ;
      RECT 2.2550 0.6800 3.0150 0.7700 ;
      RECT 2.9250 0.7700 3.0150 1.3050 ;
      RECT 2.6200 1.4700 3.2800 1.5600 ;
      RECT 2.6200 1.0500 2.7100 1.4700 ;
      RECT 3.1900 0.7700 3.2800 1.4700 ;
      RECT 3.1100 0.6800 3.2800 0.7700 ;
      RECT 3.3900 1.4700 3.9250 1.5600 ;
      RECT 3.8350 0.7700 3.9250 1.4700 ;
      RECT 3.5500 0.6800 4.2850 0.7700 ;
      RECT 4.1950 0.7700 4.2850 0.9550 ;
      RECT 4.1950 0.9550 4.3350 1.1650 ;
      RECT 1.3400 1.7700 2.1650 1.8600 ;
      RECT 2.0750 1.7400 2.1650 1.7700 ;
      RECT 1.3400 0.7500 1.4300 1.7700 ;
      RECT 2.0750 1.6500 4.8600 1.7400 ;
      RECT 1.2400 0.6600 1.4300 0.7500 ;
      RECT 4.7700 0.9500 4.8600 1.6500 ;
      RECT 4.6750 0.8600 4.8600 0.9500 ;
      RECT 4.9900 1.0500 5.3900 1.1400 ;
      RECT 4.0150 1.4200 4.5550 1.5100 ;
      RECT 4.4650 1.2100 4.5550 1.4200 ;
      RECT 4.0150 1.0250 4.1050 1.4200 ;
      RECT 4.4650 1.0400 4.6600 1.2100 ;
      RECT 4.4650 0.7700 4.5550 1.0400 ;
      RECT 4.3800 0.6800 5.0800 0.7700 ;
      RECT 4.9900 0.7700 5.0800 1.0500 ;
      RECT 2.0750 0.4800 5.9000 0.5700 ;
      RECT 5.8100 0.5700 5.9000 1.7200 ;
      RECT 3.3700 1.2700 3.7250 1.3600 ;
      RECT 3.3700 0.5700 3.4600 1.2700 ;
      RECT 2.0750 0.5700 2.1650 1.3600 ;
      RECT 2.3950 0.4100 2.5650 0.4800 ;
      RECT 6.0100 1.6500 6.5550 1.7400 ;
      RECT 6.0100 0.6000 6.5550 0.6900 ;
      RECT 2.2950 1.8300 6.1000 1.9200 ;
      RECT 6.0100 1.7400 6.1000 1.8300 ;
      RECT 6.0100 0.6900 6.1000 1.6500 ;
      RECT 3.2650 1.9200 3.4350 1.9850 ;
  END
END EDFFQN_X2M_A12TH

MACRO EDFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.7200 ;
        RECT 1.6000 0.3200 1.7700 0.3600 ;
        RECT 5.0850 0.3200 5.2550 0.3550 ;
        RECT 5.6050 0.3200 5.7750 0.3550 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.9400 6.7800 1.3900 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0606 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8350 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.105 ;
  END E

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 0.8450 5.9500 1.2900 ;
        RECT 5.3850 1.2900 6.0000 1.3900 ;
        RECT 5.3300 0.7450 6.0550 0.8450 ;
        RECT 5.3850 1.3900 5.4750 1.7200 ;
        RECT 5.9000 1.3900 6.0000 1.7250 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 0.4100 1.8950 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6900 1.4500 0.9500 1.5400 ;
      RECT 0.8500 0.6650 0.9500 1.4500 ;
      RECT 0.6750 0.5750 0.9500 0.6650 ;
      RECT 0.0500 1.7050 1.0900 1.7950 ;
      RECT 0.0500 0.6650 0.1400 1.7050 ;
      RECT 0.0500 0.5750 0.2450 0.6650 ;
      RECT 1.0600 0.5700 1.1500 1.5700 ;
      RECT 1.0600 0.4800 1.8150 0.5700 ;
      RECT 1.7250 0.5700 1.8150 1.3100 ;
      RECT 1.9250 0.5250 2.0250 1.6600 ;
      RECT 2.1600 1.4700 2.3850 1.5600 ;
      RECT 2.2950 0.7700 2.3850 1.4700 ;
      RECT 2.2950 0.6800 3.0300 0.7700 ;
      RECT 2.9400 0.7700 3.0300 0.8700 ;
      RECT 2.9400 0.8700 3.0900 1.2600 ;
      RECT 2.6600 1.4700 3.2900 1.5600 ;
      RECT 2.6600 1.0500 2.7500 1.4700 ;
      RECT 3.2000 0.7700 3.2900 1.4700 ;
      RECT 3.1200 0.6800 3.2900 0.7700 ;
      RECT 3.4000 1.4700 3.9350 1.5600 ;
      RECT 3.8450 0.7700 3.9350 1.4700 ;
      RECT 3.5600 0.6800 4.3300 0.7700 ;
      RECT 4.2400 0.7700 4.3300 0.9750 ;
      RECT 4.2400 0.9750 4.4150 1.1450 ;
      RECT 1.3750 1.7700 2.2100 1.8600 ;
      RECT 2.1200 1.7400 2.2100 1.7700 ;
      RECT 1.3750 0.7500 1.4650 1.7700 ;
      RECT 2.1200 1.6500 4.9100 1.7400 ;
      RECT 1.2800 0.6600 1.4650 0.7500 ;
      RECT 4.8200 0.9500 4.9100 1.6500 ;
      RECT 4.7250 0.8600 4.9100 0.9500 ;
      RECT 5.0650 1.0800 5.7150 1.1700 ;
      RECT 4.0250 1.4200 4.6150 1.5100 ;
      RECT 4.5250 1.2100 4.6150 1.4200 ;
      RECT 4.0250 1.0250 4.1150 1.4200 ;
      RECT 4.5250 1.0400 4.7100 1.2100 ;
      RECT 4.5250 0.7700 4.6150 1.0400 ;
      RECT 4.4300 0.6800 5.1550 0.7700 ;
      RECT 5.0650 0.7700 5.1550 1.0800 ;
      RECT 2.1150 0.4800 6.2450 0.5700 ;
      RECT 6.1550 0.5700 6.2450 1.7200 ;
      RECT 3.3800 1.2700 3.7350 1.3600 ;
      RECT 3.3800 0.5700 3.4700 1.2700 ;
      RECT 2.1150 0.5700 2.2050 1.3600 ;
      RECT 2.4350 0.4100 2.6050 0.4800 ;
      RECT 6.3550 1.6500 6.9550 1.7400 ;
      RECT 6.3550 0.6350 6.9500 0.7250 ;
      RECT 2.3350 1.8300 6.4450 1.9200 ;
      RECT 6.3550 1.7400 6.4450 1.8300 ;
      RECT 6.3550 0.7250 6.4450 1.6500 ;
      RECT 3.5200 1.9200 3.6900 1.9850 ;
  END
END EDFFQN_X3M_A12TH

MACRO EDFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.7250 ;
        RECT 1.4950 0.3200 1.7050 0.3900 ;
        RECT 5.9050 0.3200 6.0050 0.4200 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3300 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.8900 6.1700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 0.9000 5.3500 1.3150 ;
        RECT 5.2500 1.3150 5.4050 1.7050 ;
        RECT 5.2500 0.7300 5.4050 0.9000 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 4.0550 2.0200 4.2650 2.0800 ;
        RECT 4.9800 2.0200 5.1900 2.0800 ;
        RECT 5.8450 2.0200 6.0550 2.0800 ;
        RECT 2.6450 2.0150 2.8550 2.0800 ;
        RECT 1.5950 1.8500 1.6950 2.0800 ;
        RECT 0.4100 1.6400 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7950 1.3700 0.9600 1.5400 ;
      RECT 0.8600 0.7200 0.9600 1.3700 ;
      RECT 0.6750 0.6300 0.9600 0.7200 ;
      RECT 0.6150 1.6800 1.1000 1.7700 ;
      RECT 0.6150 1.5300 0.7050 1.6800 ;
      RECT 0.0500 1.4400 0.7050 1.5300 ;
      RECT 0.0500 0.7250 0.1400 1.4400 ;
      RECT 0.0500 0.5350 0.1850 0.7250 ;
      RECT 1.0600 0.5700 1.1500 1.5600 ;
      RECT 1.0600 0.4800 1.7800 0.5700 ;
      RECT 1.6900 0.5700 1.7800 1.3250 ;
      RECT 1.8550 1.4700 2.0250 1.5600 ;
      RECT 1.8950 0.6050 1.9850 1.4700 ;
      RECT 2.1400 1.4700 2.3500 1.5600 ;
      RECT 2.2600 0.7700 2.3500 1.4700 ;
      RECT 2.2600 0.6800 3.0150 0.7700 ;
      RECT 2.9250 0.7700 3.0150 1.1800 ;
      RECT 2.5600 1.4700 3.1950 1.5600 ;
      RECT 2.5600 1.1650 2.6500 1.4700 ;
      RECT 3.1050 0.7700 3.1950 1.4700 ;
      RECT 3.1050 0.6800 3.2850 0.7700 ;
      RECT 3.9600 1.4700 4.5700 1.5600 ;
      RECT 4.4800 1.2450 4.5700 1.4700 ;
      RECT 3.9600 1.1050 4.0500 1.4700 ;
      RECT 4.4800 1.0750 4.6800 1.2450 ;
      RECT 4.4800 0.9500 4.5700 1.0750 ;
      RECT 4.3950 0.8600 4.5700 0.9500 ;
      RECT 1.3200 1.6500 4.8700 1.7400 ;
      RECT 4.7200 1.3700 4.8700 1.6500 ;
      RECT 1.3200 1.3500 1.4700 1.6500 ;
      RECT 4.7800 0.9550 4.8700 1.3700 ;
      RECT 1.3800 0.7500 1.4700 1.3500 ;
      RECT 4.6800 0.8650 4.8700 0.9550 ;
      RECT 1.2600 0.6600 1.4700 0.7500 ;
      RECT 3.3050 1.4700 3.8500 1.5600 ;
      RECT 3.7600 0.7700 3.8500 1.4700 ;
      RECT 3.5550 0.6800 5.1600 0.7700 ;
      RECT 4.1950 0.7700 4.2850 1.2950 ;
      RECT 5.0700 0.7700 5.1600 1.2650 ;
      RECT 2.0800 0.4800 5.6550 0.5700 ;
      RECT 5.5650 0.5700 5.6550 1.6150 ;
      RECT 3.4550 1.2900 3.6500 1.3800 ;
      RECT 3.4550 0.9800 3.5450 1.2900 ;
      RECT 3.3750 0.8800 3.5450 0.9800 ;
      RECT 3.3750 0.5700 3.4650 0.8800 ;
      RECT 2.0800 0.5700 2.1700 1.3600 ;
      RECT 2.3350 0.4350 2.5050 0.4800 ;
      RECT 5.7750 1.6050 6.3200 1.6950 ;
      RECT 6.2300 1.4600 6.3200 1.6050 ;
      RECT 5.7750 0.6100 6.3200 0.7000 ;
      RECT 6.2300 0.7000 6.3200 0.8200 ;
      RECT 2.2500 1.8300 5.8650 1.9200 ;
      RECT 5.7750 1.6950 5.8650 1.8300 ;
      RECT 5.7750 0.7000 5.8650 1.6050 ;
  END
END EDFFQ_X0P5M_A12TH

MACRO EDFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6350 ;
        RECT 1.5250 0.3200 1.7350 0.3900 ;
        RECT 5.0050 0.3200 5.2150 0.3900 ;
        RECT 5.8950 0.3200 5.9950 0.5000 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3400 ;
    END
    ANTENNAGATEAREA 0.0702 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.8200 6.1700 1.3700 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 0.9000 5.3500 1.3150 ;
        RECT 5.2500 1.3150 5.4200 1.7050 ;
        RECT 5.2500 0.7300 5.4200 0.9000 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
        RECT 4.0550 2.0200 4.2650 2.0800 ;
        RECT 5.8400 2.0200 6.0500 2.0800 ;
        RECT 2.6450 2.0150 2.8550 2.0800 ;
        RECT 1.5400 2.0050 1.7500 2.0800 ;
        RECT 0.4100 1.6500 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7950 1.4150 0.9500 1.5850 ;
      RECT 0.8500 0.6650 0.9500 1.4150 ;
      RECT 0.7150 0.5750 0.9500 0.6650 ;
      RECT 0.6150 1.7550 1.0800 1.8450 ;
      RECT 0.6150 1.5400 0.7050 1.7550 ;
      RECT 0.0500 1.4500 0.7050 1.5400 ;
      RECT 0.0500 0.6550 0.1400 1.4500 ;
      RECT 0.0500 0.5650 0.2450 0.6550 ;
      RECT 1.0600 0.5700 1.1500 1.5650 ;
      RECT 1.0600 0.4800 1.7800 0.5700 ;
      RECT 1.6900 0.5700 1.7800 1.3250 ;
      RECT 1.8550 1.4700 2.0250 1.5600 ;
      RECT 1.8900 0.5000 1.9900 1.4700 ;
      RECT 2.1400 1.4700 2.3500 1.5600 ;
      RECT 2.2600 0.7700 2.3500 1.4700 ;
      RECT 2.2600 0.6800 3.0150 0.7700 ;
      RECT 2.9250 0.7700 3.0150 1.1800 ;
      RECT 2.5600 1.4700 3.1950 1.5600 ;
      RECT 2.5600 1.1650 2.6500 1.4700 ;
      RECT 3.1050 0.7700 3.1950 1.4700 ;
      RECT 3.1050 0.6800 3.2850 0.7700 ;
      RECT 3.9600 1.4700 4.5850 1.5600 ;
      RECT 4.4950 1.1900 4.5850 1.4700 ;
      RECT 3.9600 1.1050 4.0500 1.4700 ;
      RECT 4.4950 1.1000 4.6950 1.1900 ;
      RECT 4.4950 0.9500 4.5850 1.1000 ;
      RECT 4.4100 0.8600 4.5850 0.9500 ;
      RECT 1.3200 1.6500 4.8850 1.7400 ;
      RECT 4.7350 1.3700 4.8850 1.6500 ;
      RECT 1.3200 0.7500 1.4100 1.6500 ;
      RECT 4.7950 0.9500 4.8850 1.3700 ;
      RECT 1.2800 0.6600 1.4500 0.7500 ;
      RECT 4.6950 0.8600 4.8850 0.9500 ;
      RECT 3.3050 1.4700 3.8500 1.5600 ;
      RECT 3.7600 0.7700 3.8500 1.4700 ;
      RECT 3.5550 0.6800 5.1600 0.7700 ;
      RECT 4.2000 0.7700 4.2900 1.2950 ;
      RECT 5.0700 0.7700 5.1600 1.2450 ;
      RECT 2.0800 0.4800 5.6700 0.5700 ;
      RECT 5.5800 0.5700 5.6700 1.6100 ;
      RECT 3.3750 1.2900 3.6500 1.3800 ;
      RECT 3.3750 0.5700 3.4650 1.2900 ;
      RECT 2.0800 0.5700 2.1700 1.3550 ;
      RECT 2.3350 0.4350 2.5050 0.4800 ;
      RECT 5.7900 1.4800 6.3500 1.5700 ;
      RECT 5.7900 0.6200 6.3500 0.7100 ;
      RECT 2.2500 1.8300 5.8800 1.9200 ;
      RECT 5.7900 1.5700 5.8800 1.8300 ;
      RECT 5.7900 0.7100 5.8800 1.4800 ;
      RECT 3.2300 1.9200 3.4000 1.9650 ;
  END
END EDFFQ_X1M_A12TH

MACRO EDFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6900 ;
        RECT 1.6400 0.3200 1.8100 0.4200 ;
        RECT 4.1450 0.3200 4.5350 0.3700 ;
        RECT 5.1450 0.3200 5.3150 0.3650 ;
        RECT 5.6650 0.3200 5.8350 0.3600 ;
        RECT 6.2900 0.3200 6.3900 0.5350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0516 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.8550 6.5500 1.2800 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9500 5.7500 1.2500 ;
        RECT 5.4450 1.2500 5.7500 1.3500 ;
        RECT 5.4450 0.8500 5.7500 0.9500 ;
        RECT 5.4450 1.3500 5.5350 1.7200 ;
        RECT 5.4450 0.7100 5.5350 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 4.1050 2.0200 4.2750 2.0800 ;
        RECT 6.2550 2.0200 6.4250 2.0800 ;
        RECT 2.8400 2.0150 3.0100 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
        RECT 1.6250 1.8300 1.7450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.4850 0.9500 1.5750 ;
      RECT 0.8500 0.6650 0.9500 1.4850 ;
      RECT 0.6800 0.5750 0.9500 0.6650 ;
      RECT 0.9000 1.7550 1.0700 1.8200 ;
      RECT 0.0500 1.6650 1.0700 1.7550 ;
      RECT 0.0500 0.6550 0.1400 1.6650 ;
      RECT 0.0500 0.5650 0.2450 0.6550 ;
      RECT 1.0400 0.6350 1.1300 1.5350 ;
      RECT 1.0400 0.5450 1.8250 0.6350 ;
      RECT 1.7350 0.6350 1.8250 1.3100 ;
      RECT 1.8800 1.4700 2.0900 1.5600 ;
      RECT 1.9350 0.5300 2.0350 1.4700 ;
      RECT 2.2050 1.4700 2.3950 1.5600 ;
      RECT 2.3050 0.7700 2.3950 1.4700 ;
      RECT 2.3050 0.6800 3.0200 0.7700 ;
      RECT 2.9300 0.7700 3.0200 1.1200 ;
      RECT 2.6650 1.4700 3.2800 1.5600 ;
      RECT 2.6650 1.0350 2.7550 1.4700 ;
      RECT 3.1900 0.7700 3.2800 1.4700 ;
      RECT 3.1100 0.6800 3.2800 0.7700 ;
      RECT 4.0350 1.4200 4.6600 1.5100 ;
      RECT 4.0350 1.1050 4.1250 1.4200 ;
      RECT 4.5700 0.9500 4.6600 1.4200 ;
      RECT 4.4550 0.8600 4.6600 0.9500 ;
      RECT 1.3800 1.6500 5.0000 1.7400 ;
      RECT 4.7950 0.9500 4.8850 1.6500 ;
      RECT 1.3800 0.8150 1.4700 1.6500 ;
      RECT 4.7950 0.8600 5.0000 0.9500 ;
      RECT 1.2400 0.7250 1.4700 0.8150 ;
      RECT 5.1200 1.0550 5.5400 1.1450 ;
      RECT 3.3900 1.4700 3.9450 1.5600 ;
      RECT 3.8550 0.7700 3.9450 1.4700 ;
      RECT 3.5700 0.6800 5.2100 0.7700 ;
      RECT 4.2400 0.7700 4.3300 1.1450 ;
      RECT 5.1200 0.7700 5.2100 1.0550 ;
      RECT 4.2400 1.1450 4.4400 1.2350 ;
      RECT 2.1250 0.4800 6.0650 0.5700 ;
      RECT 5.9750 0.5700 6.0650 1.5450 ;
      RECT 3.5750 1.2900 3.7450 1.3800 ;
      RECT 3.5750 0.9700 3.6650 1.2900 ;
      RECT 3.3900 0.8800 3.6650 0.9700 ;
      RECT 3.3900 0.5700 3.4800 0.8800 ;
      RECT 2.1250 0.5700 2.2150 1.3600 ;
      RECT 2.4350 0.4100 2.6050 0.4800 ;
      RECT 6.1750 1.4800 6.7500 1.5700 ;
      RECT 6.1750 0.6300 6.7500 0.7200 ;
      RECT 2.3900 1.8300 6.2650 1.9200 ;
      RECT 6.1750 1.5700 6.2650 1.8300 ;
      RECT 6.1750 0.7200 6.2650 1.4800 ;
      RECT 3.5700 1.9200 3.7400 1.9800 ;
  END
END EDFFQ_X2M_A12TH

MACRO EDFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.0450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6900 ;
        RECT 1.6400 0.3200 1.8100 0.4200 ;
        RECT 2.8800 0.3200 2.9700 0.3600 ;
        RECT 4.1450 0.3200 4.5350 0.3700 ;
        RECT 5.1200 0.3200 5.2900 0.3650 ;
        RECT 5.6400 0.3200 5.8100 0.3600 ;
        RECT 6.5050 0.3200 6.6050 0.5350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8500 0.7500 1.2700 ;
    END
    ANTENNAGATEAREA 0.0576 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8500 0.3500 1.2700 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END E

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.9650 6.7700 1.3900 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4200 1.2500 6.0300 1.3500 ;
        RECT 5.4200 1.3500 5.5100 1.7200 ;
        RECT 5.9400 1.3500 6.0300 1.7200 ;
        RECT 5.9300 0.9500 6.0300 1.2500 ;
        RECT 5.4200 0.8500 6.0300 0.9500 ;
        RECT 5.4200 0.6900 5.5100 0.8500 ;
        RECT 5.9400 0.6900 6.0300 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.0450 2.7200 ;
        RECT 4.1050 2.0200 4.2750 2.0800 ;
        RECT 6.4700 2.0200 6.6400 2.0800 ;
        RECT 2.8400 2.0150 3.0100 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
        RECT 1.6250 1.8300 1.7450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.4850 0.9500 1.5750 ;
      RECT 0.8600 0.6650 0.9500 1.4850 ;
      RECT 0.6800 0.5750 0.9500 0.6650 ;
      RECT 0.9000 1.7550 1.0700 1.8200 ;
      RECT 0.0500 1.6650 1.0700 1.7550 ;
      RECT 0.0500 0.6550 0.1400 1.6650 ;
      RECT 0.0500 0.5650 0.2450 0.6550 ;
      RECT 1.0400 0.6350 1.1300 1.5250 ;
      RECT 1.0400 0.5450 1.8250 0.6350 ;
      RECT 1.7350 0.6350 1.8250 1.2950 ;
      RECT 1.8800 1.4700 2.0900 1.5600 ;
      RECT 1.9350 0.5300 2.0350 1.4700 ;
      RECT 2.2050 1.4700 2.4050 1.5600 ;
      RECT 2.3150 0.7800 2.4050 1.4700 ;
      RECT 2.3150 0.6900 3.0200 0.7800 ;
      RECT 2.9300 0.7800 3.0200 1.1600 ;
      RECT 2.6650 1.4700 3.2800 1.5600 ;
      RECT 2.6650 1.0350 2.7550 1.4700 ;
      RECT 3.1900 0.7700 3.2800 1.4700 ;
      RECT 3.1100 0.6800 3.2800 0.7700 ;
      RECT 4.0350 1.4200 4.6850 1.5100 ;
      RECT 4.0350 1.1050 4.1250 1.4200 ;
      RECT 4.5950 0.9500 4.6850 1.4200 ;
      RECT 4.4400 0.8600 4.6850 0.9500 ;
      RECT 1.3800 1.6500 4.9650 1.7400 ;
      RECT 4.8750 0.9500 4.9650 1.6500 ;
      RECT 1.3800 0.8150 1.4700 1.6500 ;
      RECT 4.7950 0.8600 4.9650 0.9500 ;
      RECT 1.2600 0.7250 1.4700 0.8150 ;
      RECT 5.0950 1.0550 5.7700 1.1450 ;
      RECT 3.3900 1.4700 3.9450 1.5600 ;
      RECT 3.8550 0.7700 3.9450 1.4700 ;
      RECT 3.5700 0.6800 5.1850 0.7700 ;
      RECT 4.2400 0.7700 4.3300 1.1450 ;
      RECT 5.0950 0.7700 5.1850 1.0550 ;
      RECT 4.2400 1.1450 4.4400 1.2350 ;
      RECT 2.1250 0.4800 6.2800 0.5700 ;
      RECT 6.1900 0.5700 6.2800 1.5200 ;
      RECT 3.3900 1.2900 3.7450 1.3800 ;
      RECT 3.3900 0.5700 3.4800 1.2900 ;
      RECT 2.1250 0.5700 2.2150 1.3600 ;
      RECT 2.4350 0.4100 2.6050 0.4800 ;
      RECT 2.3900 1.8300 6.9200 1.9200 ;
      RECT 6.8300 1.4800 6.9200 1.8300 ;
      RECT 6.3800 0.7550 6.9200 0.8450 ;
      RECT 6.8300 0.5850 6.9200 0.7550 ;
      RECT 6.3800 0.8450 6.4700 1.8300 ;
      RECT 3.5700 1.9200 3.7400 1.9850 ;
  END
END EDFFQ_X3M_A12TH

MACRO ENDCAPTIE2_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.4450 2.7200 ;
        RECT 0.1500 1.4500 0.2500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.4450 0.3200 ;
        RECT 0.1500 0.3200 0.2500 0.8450 ;
    END
  END VSS
END ENDCAPTIE2_A12TH

MACRO ESDFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6900 ;
        RECT 2.3850 0.3200 2.5550 0.4700 ;
        RECT 2.9250 0.3200 3.0950 0.4900 ;
        RECT 4.1250 0.3200 4.2950 0.3900 ;
        RECT 6.3700 0.3200 6.5400 0.3550 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0555 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9700 2.7600 1.3550 ;
    END
    ANTENNAGATEAREA 0.0456 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 0.9950 2.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.8200 7.5700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.9000 6.7500 1.5300 ;
        RECT 6.6500 1.5300 6.8150 1.7000 ;
        RECT 6.6500 0.7300 6.8150 0.9000 ;
    END
    ANTENNADIFFAREA 0.1304 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 5.4750 2.0200 5.6450 2.0800 ;
        RECT 7.2550 2.0200 7.4250 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
        RECT 2.4100 1.8400 2.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.4800 0.4800 7.0650 0.5700 ;
      RECT 6.9750 0.5700 7.0650 1.6250 ;
      RECT 4.8800 1.2800 5.0650 1.3700 ;
      RECT 4.8800 0.9600 4.9700 1.2800 ;
      RECT 4.7000 0.8700 4.9700 0.9600 ;
      RECT 4.7550 0.5700 4.8450 0.8700 ;
      RECT 3.4800 0.5700 3.5700 1.3600 ;
      RECT 3.7650 0.4100 3.9350 0.4800 ;
      RECT 7.1650 1.4800 7.7550 1.5700 ;
      RECT 7.1650 0.6300 7.7550 0.7200 ;
      RECT 3.7300 1.8300 7.2550 1.9200 ;
      RECT 7.1650 1.5700 7.2550 1.8300 ;
      RECT 7.1650 0.7200 7.2550 1.4800 ;
      RECT 3.7300 1.9200 3.9000 1.9650 ;
      RECT 0.7500 1.4600 0.9500 1.5500 ;
      RECT 0.8500 0.6900 0.9500 1.4600 ;
      RECT 0.7350 0.6000 0.9500 0.6900 ;
      RECT 0.7950 1.8800 1.1250 1.9700 ;
      RECT 0.7950 1.7300 0.8850 1.8800 ;
      RECT 0.0500 1.6400 0.8850 1.7300 ;
      RECT 0.0500 0.6900 0.1400 1.6400 ;
      RECT 0.0500 0.6000 0.2250 0.6900 ;
      RECT 1.0600 0.5700 1.1500 1.6750 ;
      RECT 1.0600 0.4800 1.6600 0.5700 ;
      RECT 1.5700 0.5700 1.6600 1.6600 ;
      RECT 2.0100 1.4700 2.8900 1.5600 ;
      RECT 2.0100 0.7700 2.8850 0.8600 ;
      RECT 2.0100 0.8600 2.1000 1.4700 ;
      RECT 1.8300 0.5800 3.1800 0.6700 ;
      RECT 3.0900 0.6700 3.1800 1.3250 ;
      RECT 1.8300 0.6700 1.9200 1.6600 ;
      RECT 3.2900 0.6150 3.3900 1.6200 ;
      RECT 3.5400 1.4700 3.7500 1.5600 ;
      RECT 3.6600 0.7700 3.7500 1.4700 ;
      RECT 3.6600 0.6800 4.4000 0.7700 ;
      RECT 4.3100 0.7700 4.4000 1.2750 ;
      RECT 3.9600 1.4700 4.5800 1.5600 ;
      RECT 3.9600 1.1850 4.0500 1.4700 ;
      RECT 4.4900 0.7700 4.5800 1.4700 ;
      RECT 4.4900 0.6800 4.6650 0.7700 ;
      RECT 4.7200 1.4700 5.2650 1.5600 ;
      RECT 5.1750 0.7600 5.2650 1.4700 ;
      RECT 4.9550 0.6700 5.6900 0.7600 ;
      RECT 5.6000 0.7600 5.6900 1.2750 ;
      RECT 2.0300 1.6500 2.7850 1.7400 ;
      RECT 2.6950 1.7400 2.7850 1.7650 ;
      RECT 2.6950 1.7650 3.6200 1.8550 ;
      RECT 3.5300 1.7400 3.6200 1.7650 ;
      RECT 3.5300 1.6500 6.2900 1.7400 ;
      RECT 6.1200 1.5200 6.2900 1.6500 ;
      RECT 6.2000 0.9500 6.2900 1.5200 ;
      RECT 6.0800 0.8600 6.2900 0.9500 ;
      RECT 1.3200 1.7700 2.1200 1.8600 ;
      RECT 2.0300 1.7400 2.1200 1.7700 ;
      RECT 1.3200 0.7500 1.4100 1.7700 ;
      RECT 1.2800 0.6600 1.4500 0.7500 ;
      RECT 5.3600 1.4700 5.9850 1.5600 ;
      RECT 5.8050 1.2350 5.8950 1.4700 ;
      RECT 5.3600 1.1050 5.4500 1.4700 ;
      RECT 5.8050 1.0600 6.0500 1.2350 ;
      RECT 5.8050 0.7600 5.8950 1.0600 ;
      RECT 5.8050 0.6700 6.5600 0.7600 ;
      RECT 6.4700 0.7600 6.5600 1.2450 ;
  END
END ESDFFQN_X0P5M_A12TH

MACRO ESDFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6900 ;
        RECT 2.3850 0.3200 2.5550 0.4700 ;
        RECT 6.4250 0.3200 6.5950 0.3550 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6000 0.9950 2.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 0.9950 2.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.8200 7.5700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.9000 6.7500 1.3150 ;
        RECT 6.6500 1.3150 6.8150 1.7050 ;
        RECT 6.6500 0.7300 6.8150 0.9000 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 5.4750 2.0200 5.6450 2.0800 ;
        RECT 7.2550 2.0200 7.4250 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
        RECT 2.4100 1.8400 2.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.4800 0.4800 7.0650 0.5700 ;
      RECT 6.9750 0.5700 7.0650 1.7200 ;
      RECT 4.8800 1.2800 5.0500 1.3700 ;
      RECT 4.8800 0.9600 4.9700 1.2800 ;
      RECT 4.7000 0.8700 4.9700 0.9600 ;
      RECT 4.7550 0.5700 4.8450 0.8700 ;
      RECT 3.4800 0.5700 3.5700 1.3550 ;
      RECT 3.7700 0.4100 3.9400 0.4800 ;
      RECT 7.1750 1.4800 7.7550 1.5700 ;
      RECT 7.1750 0.6300 7.7550 0.7200 ;
      RECT 3.7300 1.8300 7.2650 1.9200 ;
      RECT 7.1750 1.5700 7.2650 1.8300 ;
      RECT 7.1750 0.7200 7.2650 1.4800 ;
      RECT 3.7300 1.9200 3.9000 1.9650 ;
      RECT 4.6300 1.9200 4.8000 1.9650 ;
      RECT 0.7500 1.4600 0.9500 1.5500 ;
      RECT 0.8500 0.6650 0.9500 1.4600 ;
      RECT 0.7350 0.5750 0.9500 0.6650 ;
      RECT 0.7950 1.8800 1.1250 1.9700 ;
      RECT 0.7950 1.7300 0.8850 1.8800 ;
      RECT 0.0500 1.6400 0.8850 1.7300 ;
      RECT 0.0500 0.6550 0.1400 1.6400 ;
      RECT 0.0500 0.5650 0.2250 0.6550 ;
      RECT 1.0600 0.5700 1.1500 1.7600 ;
      RECT 1.0600 0.4800 1.6600 0.5700 ;
      RECT 1.5700 0.5700 1.6600 1.6600 ;
      RECT 2.0100 1.4700 2.8900 1.5600 ;
      RECT 2.0100 0.7700 2.8850 0.8600 ;
      RECT 2.0100 0.8600 2.1000 1.4700 ;
      RECT 1.8300 0.5800 3.1800 0.6700 ;
      RECT 3.0900 0.6700 3.1800 1.3250 ;
      RECT 1.8300 0.6700 1.9200 1.6600 ;
      RECT 3.2900 0.6850 3.3900 1.7300 ;
      RECT 3.2950 0.5150 3.3850 0.6850 ;
      RECT 3.5400 1.4700 3.7500 1.5600 ;
      RECT 3.6600 0.7700 3.7500 1.4700 ;
      RECT 3.6600 0.6800 4.4000 0.7700 ;
      RECT 4.3100 0.7700 4.4000 1.2750 ;
      RECT 3.9600 1.4700 4.5800 1.5600 ;
      RECT 3.9600 1.1850 4.0500 1.4700 ;
      RECT 4.4900 0.7700 4.5800 1.4700 ;
      RECT 4.4900 0.6800 4.6650 0.7700 ;
      RECT 4.7050 1.4700 5.2500 1.5600 ;
      RECT 5.1600 0.7600 5.2500 1.4700 ;
      RECT 4.9550 0.6700 5.6900 0.7600 ;
      RECT 5.6000 0.7600 5.6900 1.2750 ;
      RECT 2.6950 1.8300 3.6200 1.9200 ;
      RECT 2.6950 1.7400 2.7850 1.8300 ;
      RECT 3.5300 1.7400 3.6200 1.8300 ;
      RECT 2.0300 1.6500 2.7850 1.7400 ;
      RECT 3.5300 1.6500 6.2900 1.7400 ;
      RECT 6.1200 1.5200 6.2900 1.6500 ;
      RECT 6.2000 0.9500 6.2900 1.5200 ;
      RECT 6.0800 0.8600 6.2900 0.9500 ;
      RECT 2.0300 1.7400 2.1200 1.7700 ;
      RECT 1.3200 1.7700 2.1200 1.8600 ;
      RECT 1.3200 0.7500 1.4100 1.7700 ;
      RECT 1.2800 0.6600 1.4500 0.7500 ;
      RECT 5.3600 1.4700 5.9850 1.5600 ;
      RECT 5.8050 1.2350 5.8950 1.4700 ;
      RECT 5.3600 1.1050 5.4500 1.4700 ;
      RECT 5.8050 1.0600 6.0500 1.2350 ;
      RECT 5.8050 0.7600 5.8950 1.0600 ;
      RECT 5.8050 0.6700 6.5600 0.7600 ;
      RECT 6.4700 0.7600 6.5600 1.2450 ;
  END
END ESDFFQN_X1M_A12TH

MACRO ESDFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.3850 0.3200 0.4850 0.6900 ;
        RECT 2.4150 0.3200 2.5850 0.4850 ;
        RECT 3.0150 0.3200 3.1850 0.5000 ;
        RECT 4.2150 0.3200 4.3850 0.3900 ;
        RECT 5.5700 0.3200 5.7400 0.3800 ;
        RECT 6.5300 0.3200 6.7000 0.3650 ;
        RECT 7.0500 0.3200 7.2200 0.3650 ;
        RECT 7.6700 0.3200 7.7700 0.5350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 0.8000 0.7600 1.1900 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8100 0.3600 1.1900 ;
    END
    ANTENNAGATEAREA 0.1002 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9950 2.7900 1.3500 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9950 2.3900 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8500 0.9650 7.9800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0500 0.9500 7.1500 1.2500 ;
        RECT 6.8300 1.2500 7.1500 1.3500 ;
        RECT 6.8300 0.8500 7.1500 0.9500 ;
        RECT 6.8300 1.3500 6.9200 1.7200 ;
        RECT 6.8300 0.7100 6.9200 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 7.6350 2.0200 7.8050 2.0800 ;
        RECT 2.4300 1.8400 2.5300 2.0800 ;
        RECT 0.3550 1.6450 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 7.5600 1.4800 8.1450 1.5700 ;
      RECT 7.5600 0.6300 8.1450 0.7200 ;
      RECT 3.7650 1.8300 7.6500 1.9200 ;
      RECT 7.5600 1.5700 7.6500 1.8300 ;
      RECT 7.5600 0.7200 7.6500 1.4800 ;
      RECT 5.1000 1.9200 5.2700 1.9800 ;
      RECT 0.6350 0.5650 0.9500 0.6650 ;
      RECT 0.8500 0.6650 0.9500 1.3400 ;
      RECT 0.7450 1.3400 0.9500 1.5950 ;
      RECT 0.8900 1.9200 1.0600 1.9700 ;
      RECT 0.5650 1.8300 1.0600 1.9200 ;
      RECT 0.5650 1.5550 0.6550 1.8300 ;
      RECT 0.0500 1.4650 0.6550 1.5550 ;
      RECT 0.0500 0.6550 0.1400 1.4650 ;
      RECT 0.0500 0.5650 0.2250 0.6550 ;
      RECT 1.0400 0.5700 1.1300 1.6850 ;
      RECT 1.0400 0.4800 1.6800 0.5700 ;
      RECT 1.5900 0.5700 1.6800 1.6600 ;
      RECT 2.0300 1.4700 2.9100 1.5600 ;
      RECT 2.0300 0.7950 2.9750 0.8850 ;
      RECT 2.0300 0.8850 2.1200 1.4700 ;
      RECT 1.8500 0.5950 3.2000 0.6850 ;
      RECT 3.1100 0.6850 3.2000 1.1500 ;
      RECT 1.8500 0.6850 1.9400 1.6600 ;
      RECT 3.2750 1.4700 3.4450 1.5600 ;
      RECT 3.3100 0.4200 3.4100 1.4700 ;
      RECT 3.6100 1.4700 3.8100 1.5600 ;
      RECT 3.7200 0.7700 3.8100 1.4700 ;
      RECT 3.7200 0.6800 4.4400 0.7700 ;
      RECT 4.3500 0.7700 4.4400 1.1200 ;
      RECT 4.0500 1.4700 4.6800 1.5600 ;
      RECT 4.0500 1.1850 4.1400 1.4700 ;
      RECT 4.5500 0.7700 4.6400 1.4700 ;
      RECT 4.5500 0.6800 4.7250 0.7700 ;
      RECT 4.8200 1.4700 5.4500 1.5600 ;
      RECT 5.3600 0.9750 5.4500 1.4700 ;
      RECT 5.3600 0.8850 5.9000 0.9750 ;
      RECT 5.8100 0.9750 5.9000 1.0550 ;
      RECT 5.3600 0.7700 5.4500 0.8850 ;
      RECT 4.9950 0.6800 5.4500 0.7700 ;
      RECT 2.0500 1.6500 6.4400 1.7400 ;
      RECT 6.3500 0.9500 6.4400 1.6500 ;
      RECT 6.1950 0.8600 6.4400 0.9500 ;
      RECT 1.3400 1.7700 2.1400 1.8600 ;
      RECT 2.0500 1.7400 2.1400 1.7700 ;
      RECT 1.3400 0.7500 1.4300 1.7700 ;
      RECT 1.2600 0.6600 1.4300 0.7500 ;
      RECT 6.5300 1.0550 6.9400 1.1450 ;
      RECT 5.5400 1.4200 6.0850 1.5100 ;
      RECT 5.9950 1.1700 6.0850 1.4200 ;
      RECT 5.5400 1.0850 5.6300 1.4200 ;
      RECT 5.9950 1.0800 6.2000 1.1700 ;
      RECT 5.9950 0.7700 6.0850 1.0800 ;
      RECT 5.8750 0.6800 6.6200 0.7700 ;
      RECT 6.5300 0.7700 6.6200 1.0550 ;
      RECT 3.5200 0.4800 7.4450 0.5700 ;
      RECT 7.3550 0.5700 7.4450 1.7300 ;
      RECT 5.0800 1.2900 5.2500 1.3800 ;
      RECT 5.0800 0.9700 5.1700 1.2900 ;
      RECT 4.8150 0.8800 5.1700 0.9700 ;
      RECT 4.8150 0.5700 4.9050 0.8800 ;
      RECT 3.5200 0.5700 3.6100 1.3800 ;
      RECT 3.8250 0.4100 3.9950 0.4800 ;
  END
END ESDFFQN_X2M_A12TH

MACRO ESDFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.4450 0.3200 ;
        RECT 0.4150 0.3200 0.5050 0.6650 ;
        RECT 2.4200 0.3200 2.5900 0.4850 ;
        RECT 3.0300 0.3200 3.2000 0.3600 ;
        RECT 4.3000 0.3200 4.3900 0.3650 ;
        RECT 6.4850 0.3200 6.6550 0.3550 ;
        RECT 7.0050 0.3200 7.1750 0.3550 ;
        RECT 7.8700 0.3200 7.9700 0.5300 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.1002 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0100 2.7800 1.4350 ;
    END
    ANTENNAGATEAREA 0.0627 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.0100 2.3800 1.4350 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0500 1.0100 8.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 0.8450 7.4000 1.2900 ;
        RECT 6.7850 1.2900 7.4000 1.3900 ;
        RECT 6.7300 0.7450 7.4000 0.8450 ;
        RECT 6.7850 1.3900 6.8750 1.7200 ;
        RECT 7.3000 1.3900 7.4000 1.7200 ;
    END
    ANTENNADIFFAREA 0.5706 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.4450 2.7200 ;
        RECT 6.4850 2.0550 6.6550 2.0800 ;
        RECT 7.0050 2.0500 7.1750 2.0800 ;
        RECT 2.4100 2.0200 2.5800 2.0800 ;
        RECT 7.8350 2.0200 8.0050 2.0800 ;
        RECT 3.0300 1.9500 3.2000 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.5150 0.4800 7.6450 0.5700 ;
      RECT 7.5550 0.5700 7.6450 1.7200 ;
      RECT 4.9650 1.2850 5.1350 1.3750 ;
      RECT 4.9650 1.0400 5.0550 1.2850 ;
      RECT 4.7800 0.9500 5.0550 1.0400 ;
      RECT 4.7800 0.5700 4.8700 0.9500 ;
      RECT 3.5150 0.5700 3.6050 1.3600 ;
      RECT 3.8350 0.4100 4.0050 0.4800 ;
      RECT 7.7550 1.5100 8.3400 1.6000 ;
      RECT 7.7550 0.7700 8.3400 0.8600 ;
      RECT 3.7550 1.8300 7.8450 1.9200 ;
      RECT 7.7550 1.6000 7.8450 1.8300 ;
      RECT 7.7550 0.8600 7.8450 1.5100 ;
      RECT 5.0050 1.9200 5.1750 1.9800 ;
      RECT 0.7100 1.4850 0.9500 1.5750 ;
      RECT 0.8500 0.6650 0.9500 1.4850 ;
      RECT 0.6950 0.5750 0.9500 0.6650 ;
      RECT 0.7000 1.8800 1.0850 1.9700 ;
      RECT 0.7000 1.7550 0.7900 1.8800 ;
      RECT 0.0500 1.6650 0.7900 1.7550 ;
      RECT 0.0500 0.6650 0.1400 1.6650 ;
      RECT 0.0500 0.5750 0.2250 0.6650 ;
      RECT 1.0400 0.5700 1.1300 1.6850 ;
      RECT 1.0400 0.4800 1.6950 0.5700 ;
      RECT 1.6050 0.5700 1.6950 1.6600 ;
      RECT 2.0450 1.5450 2.9250 1.6350 ;
      RECT 2.0450 0.7950 2.9200 0.8850 ;
      RECT 2.0450 0.8850 2.1350 1.5450 ;
      RECT 1.8650 0.5950 3.2150 0.6850 ;
      RECT 3.1250 0.6850 3.2150 1.2450 ;
      RECT 1.8650 0.6850 1.9550 1.6600 ;
      RECT 3.3250 0.4300 3.4250 1.6600 ;
      RECT 3.5800 1.4700 3.7850 1.5600 ;
      RECT 3.6950 0.7700 3.7850 1.4700 ;
      RECT 3.6950 0.6800 4.4300 0.7700 ;
      RECT 4.3400 0.7700 4.4300 0.9250 ;
      RECT 4.3400 0.9250 4.4900 1.0950 ;
      RECT 4.0600 1.3250 4.6900 1.4150 ;
      RECT 4.0600 1.0500 4.1500 1.3250 ;
      RECT 4.6000 0.7700 4.6900 1.3250 ;
      RECT 4.5200 0.6800 4.6900 0.7700 ;
      RECT 4.7650 1.4700 5.3350 1.5600 ;
      RECT 5.2450 0.7700 5.3350 1.4700 ;
      RECT 4.9600 0.6800 5.7300 0.7700 ;
      RECT 5.6400 0.7700 5.7300 0.9750 ;
      RECT 5.6400 0.9750 5.7900 1.1450 ;
      RECT 1.3550 1.7700 3.6100 1.8600 ;
      RECT 3.5200 1.7400 3.6100 1.7700 ;
      RECT 3.5200 1.6500 6.3100 1.7400 ;
      RECT 6.2200 0.9500 6.3100 1.6500 ;
      RECT 6.1250 0.8600 6.3100 0.9500 ;
      RECT 1.3550 0.7500 1.4450 1.7700 ;
      RECT 1.2600 0.6600 1.4450 0.7500 ;
      RECT 6.4650 1.0800 7.1300 1.1700 ;
      RECT 5.4250 1.4200 6.0150 1.5100 ;
      RECT 5.9250 1.2100 6.0150 1.4200 ;
      RECT 5.4250 1.0050 5.5150 1.4200 ;
      RECT 5.9250 1.0400 6.0800 1.2100 ;
      RECT 5.9250 0.7700 6.0150 1.0400 ;
      RECT 5.8300 0.6800 6.5550 0.7700 ;
      RECT 6.4650 0.7700 6.5550 1.0800 ;
  END
END ESDFFQN_X3M_A12TH

MACRO ESDFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.7250 ;
        RECT 2.4350 0.3200 2.6050 0.4850 ;
        RECT 2.9750 0.3200 3.1450 0.4850 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8400 0.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8100 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9950 2.7900 1.3500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9950 2.3900 1.3500 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.9550 7.6000 1.3450 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.9650 6.7500 1.5150 ;
        RECT 6.6500 1.5150 6.8400 1.6850 ;
        RECT 6.6500 0.7950 6.8400 0.9650 ;
    END
    ANTENNADIFFAREA 0.124 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 5.5050 2.0200 5.6750 2.0800 ;
        RECT 2.4600 1.8400 2.5600 2.0800 ;
        RECT 0.4150 1.7300 0.5150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.7450 1.4700 5.3000 1.5600 ;
      RECT 5.2100 0.7700 5.3000 1.4700 ;
      RECT 4.9850 0.6800 6.5550 0.7700 ;
      RECT 5.6300 0.7700 5.7200 1.1050 ;
      RECT 6.4650 0.7700 6.5550 1.3850 ;
      RECT 5.6300 1.1050 5.7700 1.2750 ;
      RECT 3.5300 0.4800 7.0700 0.5700 ;
      RECT 6.9800 0.5700 7.0700 1.6150 ;
      RECT 4.8050 1.2800 5.1000 1.3700 ;
      RECT 4.8050 0.5700 4.8950 1.2800 ;
      RECT 3.5300 0.5700 3.6200 1.3600 ;
      RECT 3.8150 0.4100 3.9850 0.4800 ;
      RECT 7.1800 1.4800 7.7550 1.5700 ;
      RECT 7.1800 0.5500 7.7550 0.6400 ;
      RECT 3.7200 1.8300 7.2700 1.9200 ;
      RECT 7.1800 1.5700 7.2700 1.8300 ;
      RECT 7.1800 0.6400 7.2700 1.4800 ;
      RECT 4.5600 1.9200 4.7300 1.9350 ;
      RECT 0.8050 1.5200 0.9600 1.6900 ;
      RECT 0.8600 0.7400 0.9600 1.5200 ;
      RECT 0.7350 0.6500 0.9600 0.7400 ;
      RECT 0.6250 1.8250 1.1250 1.9150 ;
      RECT 0.6250 1.6300 0.7150 1.8250 ;
      RECT 0.0500 1.5400 0.7150 1.6300 ;
      RECT 0.0500 0.7150 0.1400 1.5400 ;
      RECT 0.0500 0.6250 0.2250 0.7150 ;
      RECT 1.0700 0.5700 1.1600 1.6850 ;
      RECT 1.0700 0.4800 1.7100 0.5700 ;
      RECT 1.6200 0.5700 1.7100 1.6600 ;
      RECT 2.0600 1.4700 2.9400 1.5600 ;
      RECT 2.0600 0.7550 2.9550 0.8450 ;
      RECT 2.0600 0.8450 2.1500 1.4700 ;
      RECT 1.8800 0.5750 3.2300 0.6650 ;
      RECT 3.1400 0.6650 3.2300 1.3250 ;
      RECT 1.8800 0.6650 1.9700 1.6600 ;
      RECT 3.3050 1.4700 3.4750 1.5600 ;
      RECT 3.3400 0.6100 3.4400 1.4700 ;
      RECT 3.6150 1.4700 3.8000 1.5600 ;
      RECT 3.7100 0.7700 3.8000 1.4700 ;
      RECT 3.7100 0.6800 4.4350 0.7700 ;
      RECT 4.3450 0.7700 4.4350 1.2750 ;
      RECT 4.0250 1.4700 4.6350 1.5600 ;
      RECT 4.0250 1.0750 4.1150 1.4700 ;
      RECT 4.5450 0.7700 4.6350 1.4700 ;
      RECT 4.5450 0.6800 4.7150 0.7700 ;
      RECT 5.4100 1.4700 6.0050 1.5600 ;
      RECT 5.9150 1.2500 6.0050 1.4700 ;
      RECT 5.4100 1.1050 5.5000 1.4700 ;
      RECT 5.9150 1.0800 6.0400 1.2500 ;
      RECT 5.9150 0.9500 6.0050 1.0800 ;
      RECT 5.8350 0.8600 6.0050 0.9500 ;
      RECT 2.0800 1.6500 6.2850 1.7400 ;
      RECT 6.1200 1.5050 6.2850 1.6500 ;
      RECT 6.1950 0.9500 6.2850 1.5050 ;
      RECT 6.1150 0.8600 6.2850 0.9500 ;
      RECT 1.3700 1.7700 2.1700 1.8600 ;
      RECT 2.0800 1.7400 2.1700 1.7700 ;
      RECT 1.3700 0.7500 1.4600 1.7700 ;
      RECT 1.2900 0.6600 1.4600 0.7500 ;
  END
END ESDFFQ_X0P5M_A12TH

MACRO ESDFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6900 ;
        RECT 2.3850 0.3200 2.5550 0.4700 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.2900 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0804 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6000 0.9950 2.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2100 0.9950 2.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4500 0.8200 7.5700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6500 0.9000 6.7500 1.3150 ;
        RECT 6.6500 1.3150 6.8150 1.7050 ;
        RECT 6.6500 0.7300 6.8150 0.9000 ;
    END
    ANTENNADIFFAREA 0.244 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 2.9450 2.0450 3.1150 2.0800 ;
        RECT 5.4750 2.0200 5.6450 2.0800 ;
        RECT 7.2550 2.0200 7.4250 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
        RECT 2.4100 1.8400 2.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.7050 1.4700 5.2500 1.5600 ;
      RECT 5.1600 0.7600 5.2500 1.4700 ;
      RECT 4.9550 0.6700 6.5600 0.7600 ;
      RECT 5.6000 0.7600 5.6900 1.2750 ;
      RECT 6.4700 0.7600 6.5600 1.2450 ;
      RECT 3.4800 0.4800 7.0650 0.5700 ;
      RECT 6.9750 0.5700 7.0650 1.7200 ;
      RECT 4.8800 1.2800 5.0500 1.3700 ;
      RECT 4.8800 0.9600 4.9700 1.2800 ;
      RECT 4.7000 0.8700 4.9700 0.9600 ;
      RECT 4.7550 0.5700 4.8450 0.8700 ;
      RECT 3.4800 0.5700 3.5700 1.3550 ;
      RECT 3.7700 0.4100 3.9400 0.4800 ;
      RECT 7.1750 1.4800 7.7550 1.5700 ;
      RECT 7.1750 0.6300 7.7550 0.7200 ;
      RECT 3.6500 1.8300 7.2650 1.9200 ;
      RECT 7.1750 1.5700 7.2650 1.8300 ;
      RECT 7.1750 0.7200 7.2650 1.4800 ;
      RECT 4.6300 1.9200 4.8000 1.9650 ;
      RECT 0.7500 1.4600 0.9500 1.5500 ;
      RECT 0.8500 0.6650 0.9500 1.4600 ;
      RECT 0.7350 0.5750 0.9500 0.6650 ;
      RECT 0.7950 1.8800 1.1250 1.9700 ;
      RECT 0.7950 1.7300 0.8850 1.8800 ;
      RECT 0.0500 1.6400 0.8850 1.7300 ;
      RECT 0.0500 0.6550 0.1400 1.6400 ;
      RECT 0.0500 0.5650 0.2250 0.6550 ;
      RECT 1.0600 0.5700 1.1500 1.7600 ;
      RECT 1.0600 0.4800 1.6600 0.5700 ;
      RECT 1.5700 0.5700 1.6600 1.6600 ;
      RECT 2.0100 1.4700 2.8900 1.5600 ;
      RECT 2.0100 0.7700 2.8850 0.8600 ;
      RECT 2.0100 0.8600 2.1000 1.4700 ;
      RECT 1.8300 0.5800 3.1800 0.6700 ;
      RECT 3.0900 0.6700 3.1800 1.3250 ;
      RECT 1.8300 0.6700 1.9200 1.6600 ;
      RECT 3.2550 1.4700 3.4250 1.5600 ;
      RECT 3.2900 0.5000 3.3900 1.4700 ;
      RECT 3.5400 1.4700 3.7500 1.5600 ;
      RECT 3.6600 0.7700 3.7500 1.4700 ;
      RECT 3.6600 0.6800 4.4000 0.7700 ;
      RECT 4.3100 0.7700 4.4000 1.2750 ;
      RECT 3.9600 1.4700 4.5800 1.5600 ;
      RECT 3.9600 1.1850 4.0500 1.4700 ;
      RECT 4.4900 0.7700 4.5800 1.4700 ;
      RECT 4.4900 0.6800 4.6650 0.7700 ;
      RECT 5.3600 1.4700 5.9850 1.5600 ;
      RECT 5.8950 1.2300 5.9850 1.4700 ;
      RECT 5.3600 1.1050 5.4500 1.4700 ;
      RECT 5.8950 1.0600 6.0550 1.2300 ;
      RECT 5.8950 0.9500 5.9850 1.0600 ;
      RECT 5.8100 0.8600 5.9850 0.9500 ;
      RECT 2.0300 1.6500 6.3100 1.7400 ;
      RECT 6.2200 0.9500 6.3100 1.6500 ;
      RECT 6.0950 0.8600 6.3100 0.9500 ;
      RECT 1.3200 1.7700 2.1200 1.8600 ;
      RECT 2.0300 1.7400 2.1200 1.7700 ;
      RECT 1.3200 0.7500 1.4100 1.7700 ;
      RECT 1.2800 0.6600 1.4500 0.7500 ;
  END
END ESDFFQ_X1M_A12TH

MACRO ESDFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.4100 0.3200 0.5100 0.6900 ;
        RECT 2.4550 0.3200 2.6250 0.4850 ;
        RECT 3.0750 0.3200 3.1750 0.4950 ;
        RECT 4.1900 0.3200 4.3600 0.3800 ;
        RECT 5.5450 0.3200 5.9350 0.3700 ;
        RECT 6.5450 0.3200 6.7150 0.3800 ;
        RECT 7.0650 0.3200 7.2350 0.3800 ;
        RECT 7.6900 0.3200 7.7900 0.5350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9950 2.8000 1.3500 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9950 2.4000 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8500 0.9650 7.9500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0500 0.9500 7.1500 1.2500 ;
        RECT 6.8450 1.2500 7.1500 1.3500 ;
        RECT 6.8450 0.8500 7.1500 0.9500 ;
        RECT 6.8450 1.3500 6.9350 1.7200 ;
        RECT 6.8450 0.7100 6.9350 0.8500 ;
    END
    ANTENNADIFFAREA 0.32 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 5.5050 2.0200 5.6750 2.0800 ;
        RECT 7.6550 2.0200 7.8250 2.0800 ;
        RECT 4.2400 2.0150 4.4100 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
        RECT 2.9800 1.8500 3.1500 2.0800 ;
        RECT 2.4700 1.8400 2.5700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 7.6400 1.4800 8.1500 1.5700 ;
      RECT 7.6400 0.6300 8.1500 0.7200 ;
      RECT 3.7900 1.8300 7.7300 1.9200 ;
      RECT 7.6400 1.5700 7.7300 1.8300 ;
      RECT 7.6400 0.7200 7.7300 1.4800 ;
      RECT 4.9700 1.9200 5.1400 1.9900 ;
      RECT 0.7150 1.4850 0.9500 1.5750 ;
      RECT 0.8500 0.6650 0.9500 1.4850 ;
      RECT 0.7000 0.5750 0.9500 0.6650 ;
      RECT 0.6800 1.8800 1.0700 1.9700 ;
      RECT 0.6800 1.7550 0.7700 1.8800 ;
      RECT 0.0500 1.6650 0.7700 1.7550 ;
      RECT 0.0500 0.6550 0.1400 1.6650 ;
      RECT 0.0500 0.5650 0.2250 0.6550 ;
      RECT 1.0400 0.5700 1.1300 1.6850 ;
      RECT 1.0400 0.4800 1.7200 0.5700 ;
      RECT 1.6300 0.5700 1.7200 1.6600 ;
      RECT 2.0700 1.4700 2.9500 1.5600 ;
      RECT 2.0700 0.7950 2.9650 0.8850 ;
      RECT 2.0700 0.8850 2.1600 1.4700 ;
      RECT 1.8900 0.5950 3.2250 0.6850 ;
      RECT 3.1350 0.6850 3.2250 1.1500 ;
      RECT 1.8900 0.6850 1.9800 1.6600 ;
      RECT 3.3000 1.4700 3.4700 1.5600 ;
      RECT 3.3350 0.5300 3.4350 1.4700 ;
      RECT 3.6250 1.4700 3.7950 1.5600 ;
      RECT 3.7050 0.7700 3.7950 1.4700 ;
      RECT 3.7050 0.6800 4.4200 0.7700 ;
      RECT 4.3300 0.7700 4.4200 1.1200 ;
      RECT 4.0650 1.4700 4.6800 1.5600 ;
      RECT 4.0650 1.0350 4.1550 1.4700 ;
      RECT 4.5900 0.7700 4.6800 1.4700 ;
      RECT 4.5100 0.6800 4.6800 0.7700 ;
      RECT 5.4350 1.4200 6.0600 1.5100 ;
      RECT 5.4350 1.0500 5.5250 1.4200 ;
      RECT 5.9700 0.9500 6.0600 1.4200 ;
      RECT 5.8550 0.8600 6.0600 0.9500 ;
      RECT 2.0900 1.6500 6.3800 1.7400 ;
      RECT 6.1950 0.9500 6.2850 1.6500 ;
      RECT 6.1950 0.8600 6.3800 0.9500 ;
      RECT 1.3800 1.7700 2.1800 1.8600 ;
      RECT 2.0900 1.7400 2.1800 1.7700 ;
      RECT 1.3800 0.7500 1.4700 1.7700 ;
      RECT 1.2600 0.6600 1.4700 0.7500 ;
      RECT 6.5200 1.0550 6.9200 1.1450 ;
      RECT 4.7900 1.4700 5.3450 1.5600 ;
      RECT 5.2550 0.7700 5.3450 1.4700 ;
      RECT 4.9700 0.6800 6.6100 0.7700 ;
      RECT 5.6400 0.7700 5.7300 1.1050 ;
      RECT 6.5200 0.7700 6.6100 1.0550 ;
      RECT 5.6400 1.1050 5.7800 1.2750 ;
      RECT 3.5250 0.4800 7.4650 0.5700 ;
      RECT 7.3750 0.5700 7.4650 1.7300 ;
      RECT 4.9750 1.2900 5.1450 1.3800 ;
      RECT 4.9750 0.9700 5.0650 1.2900 ;
      RECT 4.7900 0.8800 5.0650 0.9700 ;
      RECT 4.7900 0.5700 4.8800 0.8800 ;
      RECT 3.5250 0.5700 3.6150 1.3600 ;
      RECT 3.8350 0.4100 4.0050 0.4800 ;
  END
END ESDFFQ_X2M_A12TH

MACRO ESDFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.4450 0.3200 ;
        RECT 0.4150 0.3200 0.5050 0.6650 ;
        RECT 2.4200 0.3200 2.5900 0.4850 ;
        RECT 3.0300 0.3200 3.2000 0.3600 ;
        RECT 4.3000 0.3200 4.3900 0.3650 ;
        RECT 5.5000 0.3200 5.6700 0.3800 ;
        RECT 6.4850 0.3200 6.6550 0.3550 ;
        RECT 7.0050 0.3200 7.1750 0.3550 ;
        RECT 7.8350 0.3200 8.0050 0.6700 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8000 0.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END D

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0100 2.7800 1.4350 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.0100 2.3800 1.4350 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0500 1.0100 8.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 0.8450 7.4000 1.2900 ;
        RECT 6.7850 1.2900 7.4000 1.3900 ;
        RECT 6.7300 0.7450 7.4000 0.8450 ;
        RECT 6.7850 1.3900 6.8750 1.7300 ;
        RECT 7.3000 1.3900 7.4000 1.7300 ;
    END
    ANTENNADIFFAREA 0.5634 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.4450 2.7200 ;
        RECT 2.4100 2.0200 2.5800 2.0800 ;
        RECT 5.4950 2.0200 5.6650 2.0800 ;
        RECT 7.8350 2.0200 8.0050 2.0800 ;
        RECT 3.0300 1.9500 3.2000 2.0800 ;
        RECT 0.4100 1.8550 0.5100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.5150 0.4800 7.6450 0.5700 ;
      RECT 7.5550 0.5700 7.6450 1.7200 ;
      RECT 4.9650 1.2850 5.1350 1.3750 ;
      RECT 4.9650 1.0400 5.0550 1.2850 ;
      RECT 4.7800 0.9500 5.0550 1.0400 ;
      RECT 4.7800 0.5700 4.8700 0.9500 ;
      RECT 3.5150 0.5700 3.6050 1.3600 ;
      RECT 3.8350 0.4100 4.0050 0.4800 ;
      RECT 7.7550 1.5100 8.3400 1.6000 ;
      RECT 7.7550 0.7700 8.3400 0.8600 ;
      RECT 3.7550 1.8300 7.8450 1.9200 ;
      RECT 7.7550 1.6000 7.8450 1.8300 ;
      RECT 7.7550 0.8600 7.8450 1.5100 ;
      RECT 5.0050 1.9200 5.1750 1.9800 ;
      RECT 0.7100 1.4850 0.9500 1.5750 ;
      RECT 0.8500 0.6650 0.9500 1.4850 ;
      RECT 0.6950 0.5750 0.9500 0.6650 ;
      RECT 0.7000 1.8800 1.0850 1.9700 ;
      RECT 0.7000 1.7550 0.7900 1.8800 ;
      RECT 0.0500 1.6650 0.7900 1.7550 ;
      RECT 0.0500 0.6650 0.1400 1.6650 ;
      RECT 0.0500 0.5750 0.2250 0.6650 ;
      RECT 1.0400 0.5700 1.1300 1.6850 ;
      RECT 1.0400 0.4800 1.6950 0.5700 ;
      RECT 1.6050 0.5700 1.6950 1.6600 ;
      RECT 2.0450 1.5450 2.9250 1.6350 ;
      RECT 2.0450 0.7950 2.9200 0.8850 ;
      RECT 2.0450 0.8850 2.1350 1.5450 ;
      RECT 1.8650 0.5950 3.2150 0.6850 ;
      RECT 3.1250 0.6850 3.2150 1.2450 ;
      RECT 1.8650 0.6850 1.9550 1.6600 ;
      RECT 3.3250 0.4300 3.4250 1.6600 ;
      RECT 3.5800 1.4700 3.7850 1.5600 ;
      RECT 3.6950 0.7700 3.7850 1.4700 ;
      RECT 3.6950 0.6800 4.4300 0.7700 ;
      RECT 4.3400 0.7700 4.4300 0.9250 ;
      RECT 4.3400 0.9250 4.4900 1.0950 ;
      RECT 4.0600 1.3250 4.6900 1.4150 ;
      RECT 4.0600 1.0500 4.1500 1.3250 ;
      RECT 4.6000 0.7700 4.6900 1.3250 ;
      RECT 4.5200 0.6800 4.6900 0.7700 ;
      RECT 5.4250 1.4200 6.0150 1.5100 ;
      RECT 5.9250 1.2100 6.0150 1.4200 ;
      RECT 5.4250 1.0750 5.5150 1.4200 ;
      RECT 5.9250 1.0400 6.0800 1.2100 ;
      RECT 5.9250 0.9500 6.0150 1.0400 ;
      RECT 5.8400 0.8600 6.0150 0.9500 ;
      RECT 1.3550 1.7700 3.6100 1.8600 ;
      RECT 3.5200 1.7400 3.6100 1.7700 ;
      RECT 3.5200 1.6500 6.3100 1.7400 ;
      RECT 6.2200 0.9500 6.3100 1.6500 ;
      RECT 6.1250 0.8600 6.3100 0.9500 ;
      RECT 1.3550 0.7500 1.4450 1.7700 ;
      RECT 1.2600 0.6600 1.4450 0.7500 ;
      RECT 6.4650 1.0800 7.1300 1.1700 ;
      RECT 4.7650 1.4700 5.3350 1.5600 ;
      RECT 5.2450 0.7700 5.3350 1.4700 ;
      RECT 4.9600 0.6800 6.5550 0.7700 ;
      RECT 5.6400 0.7700 5.7300 1.1050 ;
      RECT 6.4650 0.7700 6.5550 1.0800 ;
      RECT 5.6400 1.1050 5.7900 1.2750 ;
  END
END ESDFFQ_X3M_A12TH

MACRO FILL128_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 25.6450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 25.6450 0.3200 ;
    END
  END VSS
END FILL128_A12TH

MACRO FILL16_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
    END
  END VSS
END FILL16_A12TH

MACRO FILL1_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.2450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.2450 0.3200 ;
    END
  END VSS
END FILL1_A12TH

MACRO FILL2_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.4450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.4450 0.3200 ;
    END
  END VSS
END FILL2_A12TH

MACRO FILL32_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.4450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.4450 0.3200 ;
    END
  END VSS
END FILL32_A12TH

MACRO FILL4_A12TH
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
    END
  END VSS
END FILL4_A12TH

MACRO DFFRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7600 ;
        RECT 1.8900 0.3200 2.0600 0.3900 ;
        RECT 2.7800 0.3200 2.9500 0.5250 ;
        RECT 4.7100 0.3200 4.8100 0.8550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 4.6900 2.0100 4.8600 2.0800 ;
        RECT 0.0750 1.6500 0.1750 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.0050 4.9250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0350 0.2300 1.4050 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6350 1.0300 1.7650 1.4000 ;
    END
    ANTENNAGATEAREA 0.0813 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 1.4100 4.0650 1.7100 ;
        RECT 3.9650 0.6700 4.0650 1.4100 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6900 0.4300 1.7100 ;
      RECT 0.5550 1.5250 0.7900 1.6150 ;
      RECT 0.7000 1.1300 0.7900 1.5250 ;
      RECT 0.7000 1.0400 1.5050 1.1300 ;
      RECT 1.4150 1.1300 1.5050 1.4300 ;
      RECT 0.7000 0.7300 0.7900 1.0400 ;
      RECT 1.0000 1.5700 2.0000 1.6600 ;
      RECT 1.9100 0.7500 2.0000 1.5700 ;
      RECT 1.5100 0.6600 2.0000 0.7500 ;
      RECT 1.0000 1.2400 1.0900 1.5700 ;
      RECT 3.1900 1.2000 3.4650 1.2900 ;
      RECT 3.1900 0.9150 3.2800 1.2000 ;
      RECT 2.1450 0.8250 3.2800 0.9150 ;
      RECT 2.1450 0.9150 2.2350 1.7000 ;
      RECT 3.6050 1.0550 3.8600 1.1450 ;
      RECT 2.6450 1.5500 3.6950 1.6400 ;
      RECT 3.6050 1.1450 3.6950 1.5500 ;
      RECT 2.6450 1.0250 2.7350 1.5500 ;
      RECT 3.6050 0.9300 3.6950 1.0550 ;
      RECT 3.3850 0.8400 3.6950 0.9300 ;
      RECT 3.3850 0.7050 3.4750 0.8400 ;
      RECT 3.1450 0.4800 4.5200 0.5700 ;
      RECT 4.4300 0.5700 4.5200 1.6050 ;
      RECT 2.4550 0.6250 3.2350 0.7150 ;
      RECT 3.1450 0.5700 3.2350 0.6250 ;
      RECT 0.5200 0.4800 2.5450 0.5700 ;
      RECT 2.4550 0.5700 2.5450 0.6250 ;
      RECT 0.5200 0.5700 0.6100 1.4150 ;
      RECT 0.7000 1.8200 5.1200 1.9100 ;
      RECT 5.0300 0.6650 5.1200 1.8200 ;
      RECT 1.9100 1.9100 2.0800 1.9800 ;
      RECT 2.4050 1.0250 2.4950 1.8200 ;
      RECT 0.7000 1.9100 0.8000 1.9900 ;
  END
END DFFRPQ_X2M_A12TH

MACRO DFFRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7600 ;
        RECT 1.8100 0.3200 1.9800 0.3900 ;
        RECT 2.8600 0.3200 3.0300 0.5250 ;
        RECT 5.1100 0.3200 5.2100 0.8550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 5.0900 2.0100 5.2600 2.0800 ;
        RECT 0.0750 1.6500 0.1750 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 1.0050 5.3250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0350 0.2300 1.4050 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6350 0.8400 1.7650 1.2250 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0550 1.4500 4.6750 1.5500 ;
        RECT 4.0550 1.5500 4.1550 1.7100 ;
        RECT 4.5750 1.5500 4.6750 1.7100 ;
        RECT 4.0550 1.2900 4.1550 1.4500 ;
        RECT 4.5750 0.9000 4.6750 1.4500 ;
        RECT 4.0000 0.8000 4.6750 0.9000 ;
        RECT 4.5750 0.6850 4.6750 0.8000 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6900 0.4300 1.8600 ;
      RECT 0.5550 1.5250 0.7900 1.6150 ;
      RECT 0.7000 0.9300 0.7900 1.5250 ;
      RECT 0.7000 0.8400 1.5050 0.9300 ;
      RECT 1.4150 0.9300 1.5050 1.2350 ;
      RECT 0.7000 0.7300 0.7900 0.8400 ;
      RECT 1.0100 1.5700 2.1900 1.6600 ;
      RECT 2.1000 0.7500 2.1900 1.5700 ;
      RECT 1.5100 0.6600 2.1900 0.7500 ;
      RECT 1.0100 1.2100 1.1000 1.5700 ;
      RECT 3.2700 1.0850 3.6650 1.1750 ;
      RECT 3.2700 0.9150 3.3600 1.0850 ;
      RECT 2.2800 0.8250 3.3600 0.9150 ;
      RECT 2.2800 0.9150 2.3700 1.7000 ;
      RECT 3.8100 1.0550 4.4150 1.1450 ;
      RECT 2.7250 1.5500 3.9000 1.6400 ;
      RECT 3.8100 1.1450 3.9000 1.5500 ;
      RECT 2.7250 1.0150 2.8150 1.5500 ;
      RECT 3.8100 0.9300 3.9000 1.0550 ;
      RECT 3.4800 0.8400 3.9000 0.9300 ;
      RECT 3.4800 0.7050 3.5700 0.8400 ;
      RECT 3.2250 0.4800 4.9200 0.5700 ;
      RECT 4.8300 0.5700 4.9200 1.7250 ;
      RECT 2.6300 0.6250 3.3150 0.7150 ;
      RECT 3.2250 0.5700 3.3150 0.6250 ;
      RECT 0.5200 0.4800 2.7200 0.5700 ;
      RECT 2.6300 0.5700 2.7200 0.6250 ;
      RECT 0.5200 0.5700 0.6100 1.4150 ;
      RECT 0.7500 1.8200 5.5200 1.9100 ;
      RECT 5.4300 0.6650 5.5200 1.8200 ;
      RECT 2.0050 1.9100 2.1750 1.9900 ;
      RECT 2.4850 1.0150 2.5750 1.8200 ;
      RECT 0.7500 1.9100 0.8500 1.9900 ;
  END
END DFFRPQ_X3M_A12TH

MACRO DFFRPQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6750 ;
        RECT 1.8100 0.3200 1.9800 0.3900 ;
        RECT 2.8600 0.3200 3.0300 0.5250 ;
        RECT 5.3100 0.3200 5.4100 0.8550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 5.2900 2.0100 5.4600 2.0800 ;
        RECT 0.0750 1.6500 0.1750 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 1.0050 5.5250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0426 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2050 0.2300 1.3900 ;
        RECT 0.1350 1.0000 0.2300 1.2050 ;
    END
    ANTENNAGATEAREA 0.0882 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6350 0.8400 1.7650 1.2250 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0400 1.4500 4.6600 1.5500 ;
        RECT 4.0400 1.5500 4.1400 1.7100 ;
        RECT 4.5600 1.5500 4.6600 1.7100 ;
        RECT 4.0400 1.2900 4.1400 1.4500 ;
        RECT 4.5600 0.9000 4.6600 1.4500 ;
        RECT 3.9850 0.8000 4.6600 0.9000 ;
        RECT 4.5600 0.6850 4.6600 0.8000 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6900 0.4300 1.8600 ;
      RECT 0.5400 1.5250 0.7900 1.6150 ;
      RECT 0.7000 0.9300 0.7900 1.5250 ;
      RECT 0.7000 0.8400 1.5050 0.9300 ;
      RECT 1.4150 0.9300 1.5050 1.2350 ;
      RECT 0.7000 0.7300 0.7900 0.8400 ;
      RECT 1.0100 1.5700 2.1900 1.6600 ;
      RECT 2.1000 0.7500 2.1900 1.5700 ;
      RECT 1.5100 0.6600 2.1900 0.7500 ;
      RECT 1.0100 1.2100 1.1000 1.5700 ;
      RECT 3.2700 1.0850 3.6150 1.1750 ;
      RECT 3.2700 0.9150 3.3600 1.0850 ;
      RECT 2.2800 0.8250 3.3600 0.9150 ;
      RECT 2.2800 0.9150 2.3700 1.7000 ;
      RECT 3.7950 1.0550 4.4000 1.1450 ;
      RECT 2.7250 1.5500 3.8850 1.6400 ;
      RECT 3.7950 1.1450 3.8850 1.5500 ;
      RECT 2.7250 1.0150 2.8150 1.5500 ;
      RECT 3.7950 0.9300 3.8850 1.0550 ;
      RECT 3.4650 0.8400 3.8850 0.9300 ;
      RECT 3.4650 0.7050 3.5550 0.8400 ;
      RECT 3.2250 0.4800 5.1200 0.5700 ;
      RECT 5.0300 0.5700 5.1200 1.7200 ;
      RECT 2.6300 0.6250 3.3150 0.7150 ;
      RECT 3.2250 0.5700 3.3150 0.6250 ;
      RECT 0.5200 0.4800 2.7200 0.5700 ;
      RECT 2.6300 0.5700 2.7200 0.6250 ;
      RECT 0.5200 0.5700 0.6100 1.3900 ;
      RECT 0.7500 1.8200 5.7200 1.9100 ;
      RECT 5.6300 0.6650 5.7200 1.8200 ;
      RECT 2.0050 1.9100 2.1750 1.9900 ;
      RECT 2.4850 1.0150 2.5750 1.8200 ;
      RECT 0.7500 1.9100 0.8500 1.9900 ;
  END
END DFFRPQ_X4M_A12TH

MACRO DFFSQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1800 0.9000 ;
        RECT 4.2950 0.3200 4.4650 0.6700 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 1.0050 4.5500 1.4250 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1500 0.1500 1.3900 ;
        RECT 0.0500 1.0500 0.2600 1.1500 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7850 1.2900 3.9500 1.7000 ;
        RECT 3.8500 0.9400 3.9500 1.2900 ;
        RECT 3.7450 0.8400 3.9500 0.9400 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.1000 1.8250 1.3150 ;
        RECT 1.6500 1.3150 1.7500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.0900 1.5000 0.1800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.6000 1.3050 3.3150 1.3950 ;
      RECT 2.6000 1.1600 2.6900 1.3050 ;
      RECT 3.0650 0.9500 3.1550 1.3050 ;
      RECT 3.0650 0.8600 3.3300 0.9500 ;
      RECT 2.1550 1.5700 3.5050 1.6600 ;
      RECT 3.4150 1.1700 3.5050 1.5700 ;
      RECT 2.1550 0.7100 2.2450 1.5700 ;
      RECT 3.3300 1.0700 3.7100 1.1700 ;
      RECT 0.5600 0.5200 4.1300 0.6100 ;
      RECT 4.0400 0.6100 4.1300 1.7050 ;
      RECT 2.3550 0.6100 2.4450 1.4750 ;
      RECT 0.5300 1.2450 0.6500 1.4150 ;
      RECT 0.5600 0.6100 0.6500 1.2450 ;
      RECT 0.6550 1.8250 4.7500 1.9150 ;
      RECT 4.6100 1.5200 4.7500 1.8250 ;
      RECT 4.6500 0.8900 4.7500 1.5200 ;
      RECT 4.2200 0.8000 4.7500 0.8900 ;
      RECT 4.6250 0.5100 4.7500 0.8000 ;
      RECT 0.3500 0.6900 0.4400 1.6600 ;
      RECT 0.5500 1.5250 0.8300 1.6150 ;
      RECT 0.7400 0.8550 0.8300 1.5250 ;
      RECT 0.7400 0.7650 1.4950 0.8550 ;
      RECT 1.4050 0.8550 1.4950 1.3000 ;
      RECT 1.3500 1.6100 2.0450 1.7100 ;
      RECT 1.9450 0.8550 2.0450 1.6100 ;
      RECT 1.7950 0.7550 2.0450 0.8550 ;
      RECT 1.3500 1.5900 1.4500 1.6100 ;
      RECT 1.0200 1.4900 1.4500 1.5900 ;
      RECT 1.0200 1.1000 1.1200 1.4900 ;
  END
END DFFSQN_X0P5M_A12TH

MACRO DFFSQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8900 ;
        RECT 3.2200 0.3200 3.5900 0.4000 ;
        RECT 4.2950 0.3200 4.4650 0.7300 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.8750 4.5500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1500 0.1500 1.3900 ;
        RECT 0.0500 1.0500 0.2500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7800 1.2900 3.9500 1.7000 ;
        RECT 3.8500 0.9450 3.9500 1.2900 ;
        RECT 3.7150 0.8450 3.9500 0.9450 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9800 1.7500 1.2550 ;
        RECT 1.6500 1.2550 1.8600 1.3450 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 1.5850 2.0000 1.8050 2.0800 ;
        RECT 0.0800 1.5000 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0100 1.6100 2.0400 1.7000 ;
      RECT 1.9500 0.8450 2.0400 1.6100 ;
      RECT 1.7450 0.7550 2.0400 0.8450 ;
      RECT 1.0100 1.1000 1.1000 1.6100 ;
      RECT 2.6200 1.3050 3.3350 1.3950 ;
      RECT 2.6200 1.1850 2.7100 1.3050 ;
      RECT 3.1200 0.9500 3.2100 1.3050 ;
      RECT 3.1200 0.8600 3.3550 0.9500 ;
      RECT 3.3300 1.0700 3.7400 1.1700 ;
      RECT 2.1350 1.5750 3.5200 1.6650 ;
      RECT 3.4300 1.1700 3.5200 1.5750 ;
      RECT 2.1350 0.7550 2.2250 1.5750 ;
      RECT 0.5400 0.6050 0.6300 1.4100 ;
      RECT 0.5400 0.5150 1.8800 0.5200 ;
      RECT 0.5400 0.5200 4.1300 0.6050 ;
      RECT 1.7400 0.6050 4.1300 0.6100 ;
      RECT 2.3400 0.6100 2.4300 1.4450 ;
      RECT 4.0400 0.6100 4.1300 1.7000 ;
      RECT 2.2700 0.5200 2.4800 0.6050 ;
      RECT 2.2700 0.6050 2.4800 0.6100 ;
      RECT 2.2700 0.4100 2.4800 0.5200 ;
      RECT 0.7300 1.8100 4.7500 1.9100 ;
      RECT 4.6300 1.5900 4.7500 1.8100 ;
      RECT 4.2300 1.5000 4.7500 1.5900 ;
      RECT 4.6500 0.7700 4.7500 1.5000 ;
      RECT 4.5850 0.6000 4.7500 0.7700 ;
      RECT 4.2300 1.1800 4.3200 1.5000 ;
      RECT 2.3750 1.9100 2.5850 1.9900 ;
      RECT 0.7300 1.9100 0.9000 1.9900 ;
      RECT 0.3400 0.4800 0.4300 1.8500 ;
      RECT 0.5400 1.5050 0.8350 1.5950 ;
      RECT 0.7450 0.8500 0.8350 1.5050 ;
      RECT 0.7450 0.7600 1.5000 0.8500 ;
      RECT 1.4100 0.8500 1.5000 1.3000 ;
  END
END DFFSQN_X1M_A12TH

MACRO DFFSQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 3.9950 0.3200 4.6300 0.3950 ;
        RECT 0.0800 0.3200 0.1700 0.6950 ;
        RECT 1.0200 0.3200 1.3900 0.3950 ;
        RECT 3.2150 0.3200 3.5850 0.3950 ;
        RECT 4.5300 0.3950 4.6300 0.8550 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.9650 4.7500 1.4050 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1500 0.1500 1.3900 ;
        RECT 0.0500 1.0500 0.2500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7700 1.2500 4.1500 1.3500 ;
        RECT 3.7700 1.3500 3.8700 1.7000 ;
        RECT 4.0500 0.9050 4.1500 1.2500 ;
        RECT 3.7100 0.8050 4.1500 0.9050 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9800 1.7900 1.3450 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0800 1.6900 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.4350 0.4300 1.8900 ;
      RECT 0.5400 1.5050 0.8350 1.5950 ;
      RECT 0.7450 0.8500 0.8350 1.5050 ;
      RECT 0.7450 0.7600 1.5000 0.8500 ;
      RECT 1.4100 0.8500 1.5000 1.2600 ;
      RECT 1.0100 1.6100 1.9900 1.7000 ;
      RECT 1.9000 0.8200 1.9900 1.6100 ;
      RECT 1.7450 0.7300 1.9900 0.8200 ;
      RECT 1.0100 1.1000 1.1000 1.6100 ;
      RECT 2.6150 1.3050 3.3350 1.3950 ;
      RECT 2.6150 1.2000 2.7050 1.3050 ;
      RECT 3.1150 0.9450 3.2050 1.3050 ;
      RECT 3.1150 0.8550 3.3550 0.9450 ;
      RECT 3.4250 1.0700 3.8400 1.1600 ;
      RECT 2.0800 1.5700 3.5150 1.6600 ;
      RECT 2.0800 1.4900 2.3800 1.5700 ;
      RECT 3.4250 1.1600 3.5150 1.5700 ;
      RECT 2.0800 0.7550 2.1700 1.4900 ;
      RECT 1.7400 0.6050 4.3300 0.6100 ;
      RECT 4.2400 0.6100 4.3300 1.6200 ;
      RECT 0.5400 0.5200 4.3300 0.6050 ;
      RECT 2.3800 1.2300 2.4750 1.4000 ;
      RECT 2.3850 0.6100 2.4750 1.2300 ;
      RECT 0.5400 0.5150 1.8800 0.5200 ;
      RECT 2.3400 0.4200 2.5500 0.5200 ;
      RECT 0.5400 0.6050 0.6300 1.4100 ;
      RECT 0.7300 1.8200 4.9550 1.9200 ;
      RECT 4.8000 1.5200 4.9550 1.8200 ;
      RECT 4.8550 0.8500 4.9550 1.5200 ;
      RECT 4.7850 0.6800 4.9550 0.8500 ;
      RECT 2.4050 1.9200 2.6150 1.9900 ;
      RECT 0.7300 1.9200 0.9000 1.9900 ;
  END
END DFFSQN_X2M_A12TH

MACRO DFFSQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6850 ;
        RECT 3.2150 0.3200 3.5850 0.3950 ;
        RECT 3.9750 0.3200 4.1850 0.4100 ;
        RECT 4.9000 0.3200 5.0000 0.7650 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0400 0.8600 5.1500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1500 0.1500 1.3900 ;
        RECT 0.0500 1.0500 0.2500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7700 1.2500 4.3850 1.3500 ;
        RECT 3.7700 1.3500 3.8700 1.7000 ;
        RECT 4.2950 1.3500 4.3850 1.7000 ;
        RECT 4.2500 0.8800 4.3500 1.2500 ;
        RECT 3.7100 0.8700 4.3500 0.8800 ;
        RECT 3.7100 0.7800 4.4450 0.8700 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END QN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9800 1.7900 1.3450 ;
    END
    ANTENNAGATEAREA 0.1212 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 0.0800 1.7000 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.4350 0.4300 1.8900 ;
      RECT 0.5400 1.5050 0.8350 1.5950 ;
      RECT 0.7450 0.8500 0.8350 1.5050 ;
      RECT 0.7450 0.7600 1.5150 0.8500 ;
      RECT 1.4250 0.8500 1.5150 1.2350 ;
      RECT 1.3550 1.6100 1.9900 1.7000 ;
      RECT 1.9000 0.8200 1.9900 1.6100 ;
      RECT 1.7450 0.7300 1.9900 0.8200 ;
      RECT 1.3550 1.4200 1.4450 1.6100 ;
      RECT 1.0100 1.3300 1.4450 1.4200 ;
      RECT 1.0100 1.1000 1.1000 1.3300 ;
      RECT 2.6150 1.3050 3.3350 1.3950 ;
      RECT 2.6150 0.9450 2.7050 1.3050 ;
      RECT 2.6150 0.8550 3.3550 0.9450 ;
      RECT 3.4250 1.0700 3.8400 1.1600 ;
      RECT 2.0800 1.5700 3.5150 1.6600 ;
      RECT 2.0800 1.4900 2.3800 1.5700 ;
      RECT 3.4250 1.1600 3.5150 1.5700 ;
      RECT 2.0800 0.7550 2.1700 1.4900 ;
      RECT 1.7400 0.6050 4.7000 0.6100 ;
      RECT 4.6100 0.6100 4.7000 1.7300 ;
      RECT 0.5400 0.5200 4.7000 0.6050 ;
      RECT 2.3800 1.2300 2.4750 1.4000 ;
      RECT 2.3850 0.6100 2.4750 1.2300 ;
      RECT 0.5400 0.5150 1.8800 0.5200 ;
      RECT 2.3400 0.4200 2.5500 0.5200 ;
      RECT 0.5400 0.6050 0.6300 1.4100 ;
      RECT 0.7100 1.8200 5.3400 1.9200 ;
      RECT 5.1750 1.3600 5.3400 1.8200 ;
      RECT 5.2400 0.7500 5.3400 1.3600 ;
      RECT 5.1750 0.5800 5.3400 0.7500 ;
      RECT 2.4050 1.9200 2.6150 1.9900 ;
      RECT 0.7100 1.9200 0.9200 1.9900 ;
  END
END DFFSQN_X3M_A12TH

MACRO DFFSQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.8450 ;
        RECT 1.3450 0.3200 1.5150 0.7400 ;
        RECT 4.4650 0.3200 4.5650 0.6600 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4450 1.0000 4.6900 1.1100 ;
        RECT 4.4450 1.1100 4.5550 1.4050 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0350 0.1700 1.3900 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8400 0.6900 3.9600 1.6700 ;
    END
    ANTENNADIFFAREA 0.134925 ;
  END Q

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.2300 1.8300 1.4000 ;
        RECT 1.6500 1.0250 1.7500 1.2300 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 3.5150 1.9700 3.7250 2.0800 ;
        RECT 4.3900 1.9700 4.6000 2.0800 ;
        RECT 0.0950 1.5000 0.1850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 0.6250 0.4450 1.6450 ;
      RECT 0.7650 1.0150 1.5000 1.1050 ;
      RECT 1.4100 1.1050 1.5000 1.3050 ;
      RECT 0.5550 1.5100 0.8550 1.6000 ;
      RECT 0.7650 1.1050 0.8550 1.5100 ;
      RECT 0.7650 0.6600 0.8550 1.0150 ;
      RECT 1.0750 1.5800 2.0450 1.6700 ;
      RECT 1.9550 0.9800 2.0450 1.5800 ;
      RECT 1.8600 0.8900 2.0450 0.9800 ;
      RECT 1.8600 0.6600 1.9500 0.8900 ;
      RECT 1.0750 1.1950 1.1650 1.5800 ;
      RECT 2.1650 1.5400 3.1950 1.6300 ;
      RECT 3.1050 1.1300 3.1950 1.5400 ;
      RECT 2.1650 0.6600 2.2550 1.5400 ;
      RECT 3.1050 1.0400 3.5250 1.1300 ;
      RECT 3.2900 1.3750 3.3800 1.5000 ;
      RECT 3.2900 1.2850 3.7450 1.3750 ;
      RECT 3.6550 0.8450 3.7450 1.2850 ;
      RECT 2.6050 0.7550 3.7450 0.8450 ;
      RECT 2.6050 0.8450 2.6950 1.3950 ;
      RECT 1.6250 0.4800 4.2250 0.5700 ;
      RECT 4.1350 0.5700 4.2250 1.4800 ;
      RECT 1.1450 0.8300 1.7150 0.9200 ;
      RECT 1.6250 0.5700 1.7150 0.8300 ;
      RECT 2.3750 0.5700 2.4650 1.4050 ;
      RECT 0.5400 0.5700 0.6300 1.3850 ;
      RECT 0.5400 0.4800 1.2350 0.5700 ;
      RECT 1.1450 0.5700 1.2350 0.8300 ;
      RECT 0.6600 1.7900 4.8800 1.8800 ;
      RECT 4.7900 0.8500 4.8800 1.7900 ;
      RECT 4.3250 0.7600 4.8800 0.8500 ;
      RECT 4.7900 0.4600 4.8800 0.7600 ;
  END
END DFFSQ_X0P5M_A12TH

MACRO DFFSQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8050 ;
        RECT 1.3600 0.3200 1.5300 0.7150 ;
        RECT 2.9350 0.3200 3.1450 0.5350 ;
        RECT 3.6350 0.3200 3.7250 0.4600 ;
        RECT 4.4650 0.3200 4.5550 0.9250 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.1400 1.8350 1.3100 ;
        RECT 1.6500 1.3100 1.7600 1.4650 ;
        RECT 1.6500 1.0500 1.7600 1.1400 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 1.1650 4.5500 1.4950 ;
        RECT 4.4500 1.0750 4.6750 1.1650 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.7850 3.9900 1.6700 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0800 1.7100 0.1700 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 0.7250 0.4300 1.7750 ;
      RECT 0.5400 1.6100 0.8500 1.7000 ;
      RECT 0.7600 1.2000 0.8500 1.6100 ;
      RECT 0.7600 1.1100 1.5400 1.2000 ;
      RECT 0.7600 0.7450 0.8500 1.1100 ;
      RECT 1.0550 1.6350 2.0500 1.7250 ;
      RECT 1.9600 0.8750 2.0500 1.6350 ;
      RECT 1.8300 0.7850 2.0500 0.8750 ;
      RECT 1.0550 1.2900 1.1450 1.6350 ;
      RECT 2.1450 1.6500 3.1850 1.7400 ;
      RECT 3.0950 1.1700 3.1850 1.6500 ;
      RECT 2.1450 0.7250 2.2350 1.6500 ;
      RECT 3.0950 1.0800 3.5100 1.1700 ;
      RECT 3.3050 1.3800 3.3950 1.7200 ;
      RECT 3.3050 1.2900 3.7300 1.3800 ;
      RECT 3.6400 0.9350 3.7300 1.2900 ;
      RECT 2.5900 0.8450 3.7300 0.9350 ;
      RECT 2.5900 0.9350 2.6800 1.5550 ;
      RECT 2.3600 0.6350 4.2500 0.6600 ;
      RECT 4.1600 0.6600 4.2500 1.5000 ;
      RECT 3.3850 0.5700 4.2500 0.6350 ;
      RECT 2.3600 0.6600 3.4750 0.7250 ;
      RECT 1.1500 0.6050 1.2400 0.8100 ;
      RECT 0.5250 0.5150 1.2400 0.6050 ;
      RECT 0.5250 0.6050 0.6150 1.4650 ;
      RECT 1.1500 0.8100 1.7400 0.9000 ;
      RECT 1.6500 0.5700 1.7400 0.8100 ;
      RECT 1.6500 0.4800 2.4950 0.5700 ;
      RECT 2.3600 0.5700 2.4950 0.6350 ;
      RECT 2.3600 0.7250 2.4500 1.5450 ;
      RECT 0.6700 1.8300 4.8900 1.9200 ;
      RECT 4.8000 0.7150 4.8900 1.8300 ;
      RECT 2.0150 1.9200 2.2250 1.9850 ;
  END
END DFFSQ_X1M_A12TH

MACRO DFFSQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9150 ;
        RECT 1.3300 0.3200 1.5000 0.6500 ;
        RECT 2.9350 0.3200 3.1450 0.4700 ;
        RECT 3.5950 0.3200 3.7650 0.5550 ;
        RECT 4.1150 0.3200 4.2850 0.5550 ;
        RECT 4.7200 0.3200 4.8200 0.7500 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 0.0800 1.5800 0.1700 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.9500 4.1500 1.2800 ;
        RECT 3.8950 1.2800 4.1500 1.3800 ;
        RECT 3.8500 0.8500 4.1500 0.9500 ;
        RECT 3.8950 1.3800 3.9850 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.1300 4.9000 1.3000 ;
        RECT 4.6500 1.3000 4.7500 1.5600 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END CK

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.2200 1.7500 1.4450 ;
        RECT 1.6500 1.0500 1.8050 1.2200 ;
    END
    ANTENNAGATEAREA 0.075 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0600 0.1800 1.4300 ;
    END
    ANTENNAGATEAREA 0.0474 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 0.5550 0.4300 1.9600 ;
      RECT 0.5400 1.6250 0.8150 1.7150 ;
      RECT 0.7250 1.2000 0.8150 1.6250 ;
      RECT 0.7250 1.1100 1.5200 1.2000 ;
      RECT 0.7250 0.7450 0.8150 1.1100 ;
      RECT 1.0200 1.6300 2.0050 1.7300 ;
      RECT 1.9050 0.8800 2.0050 1.6300 ;
      RECT 1.7800 0.7800 2.0050 0.8800 ;
      RECT 1.0200 1.2900 1.1200 1.6300 ;
      RECT 2.1250 1.6500 3.1850 1.7400 ;
      RECT 3.0950 1.1700 3.1850 1.6500 ;
      RECT 2.1250 0.7250 2.2150 1.6500 ;
      RECT 3.0950 1.0800 3.5100 1.1700 ;
      RECT 3.6650 1.0800 3.9550 1.1700 ;
      RECT 3.2950 1.3800 3.3850 1.7200 ;
      RECT 3.2950 1.2900 3.7550 1.3800 ;
      RECT 3.6650 1.1700 3.7550 1.2900 ;
      RECT 3.6650 0.9350 3.7550 1.0800 ;
      RECT 2.5900 0.8450 3.7550 0.9350 ;
      RECT 2.5900 0.9350 2.6800 1.5400 ;
      RECT 2.3600 0.6450 4.5100 0.7350 ;
      RECT 4.4200 0.7350 4.5100 1.7400 ;
      RECT 1.1200 0.6050 1.2100 0.7500 ;
      RECT 0.5250 0.5150 1.2100 0.6050 ;
      RECT 0.5250 0.6050 0.6150 1.5100 ;
      RECT 1.1200 0.7500 1.6900 0.8400 ;
      RECT 1.6000 0.5700 1.6900 0.7500 ;
      RECT 1.6000 0.4800 2.4500 0.5700 ;
      RECT 2.3600 0.5700 2.4500 0.6450 ;
      RECT 2.0000 0.4100 2.1700 0.4800 ;
      RECT 2.3600 0.7350 2.4500 1.5500 ;
      RECT 0.6700 1.8300 5.1050 1.9200 ;
      RECT 5.0150 1.0000 5.1050 1.8300 ;
      RECT 4.6000 0.9100 5.1050 1.0000 ;
      RECT 5.0150 0.6100 5.1050 0.9100 ;
      RECT 0.6700 1.9200 0.8800 1.9900 ;
      RECT 2.0050 1.9200 2.2150 1.9850 ;
  END
END DFFSQ_X2M_A12TH

MACRO DFFSQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.9300 ;
        RECT 1.3700 0.3200 1.4600 0.5600 ;
        RECT 3.5600 0.3200 3.7300 0.5200 ;
        RECT 4.0800 0.3200 4.2500 0.5100 ;
        RECT 4.9500 0.3200 5.0500 0.6750 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6450 1.0300 1.8150 1.4150 ;
    END
    ANTENNAGATEAREA 0.0882 ;
  END SN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8550 1.2500 4.5500 1.3500 ;
        RECT 3.8550 1.3500 3.9550 1.6900 ;
        RECT 4.3800 1.3500 4.4700 1.6700 ;
        RECT 4.4500 0.9100 4.5500 1.2500 ;
        RECT 3.8200 0.8100 4.5500 0.9100 ;
    END
    ANTENNADIFFAREA 0.595725 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.2350 4.9500 1.6000 ;
        RECT 4.8500 1.1350 5.1350 1.2350 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 1.5700 2.0050 1.7800 2.0800 ;
        RECT 0.0950 1.5200 0.1850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 0.5200 0.4450 1.8800 ;
      RECT 0.5650 1.4950 0.8450 1.5850 ;
      RECT 0.7550 0.9200 0.8450 1.4950 ;
      RECT 0.7550 0.8300 1.5250 0.9200 ;
      RECT 1.4350 0.9200 1.5250 1.2400 ;
      RECT 1.0900 1.5800 2.0350 1.6700 ;
      RECT 1.9450 0.8000 2.0350 1.5800 ;
      RECT 1.7700 0.7100 2.0350 0.8000 ;
      RECT 1.0900 1.1900 1.1800 1.5800 ;
      RECT 2.1550 1.4700 3.2400 1.5600 ;
      RECT 3.1500 1.1600 3.2400 1.4700 ;
      RECT 2.1550 0.7850 2.2450 1.4700 ;
      RECT 3.1500 1.0600 3.5450 1.1600 ;
      RECT 3.6400 1.0550 4.2700 1.1450 ;
      RECT 3.3400 1.3750 3.4300 1.7050 ;
      RECT 3.3400 1.2750 3.7300 1.3750 ;
      RECT 3.6400 1.1450 3.7300 1.2750 ;
      RECT 3.6400 0.8900 3.7300 1.0550 ;
      RECT 2.6500 0.8000 3.7300 0.8900 ;
      RECT 2.6500 0.8900 2.7400 1.3650 ;
      RECT 2.3900 0.6100 4.7350 0.7000 ;
      RECT 4.6450 0.7000 4.7350 1.7350 ;
      RECT 0.5450 0.7400 0.6350 1.3850 ;
      RECT 0.8350 0.5950 1.0450 0.6500 ;
      RECT 0.5450 0.6500 1.6600 0.7400 ;
      RECT 1.5700 0.5700 1.6600 0.6500 ;
      RECT 1.5700 0.4800 2.4800 0.5700 ;
      RECT 2.3900 0.5700 2.4800 0.6100 ;
      RECT 2.3900 0.7000 2.4800 1.3800 ;
      RECT 0.7650 1.8250 5.3200 1.9150 ;
      RECT 5.2300 0.9700 5.3200 1.8250 ;
      RECT 4.8250 0.8800 5.3200 0.9700 ;
      RECT 5.2300 0.5850 5.3200 0.8800 ;
      RECT 2.2950 1.9150 2.5050 1.9900 ;
      RECT 0.7650 1.9150 0.9350 1.9800 ;
  END
END DFFSQ_X3M_A12TH

MACRO DFFSQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.0900 0.3200 0.1800 0.8350 ;
        RECT 1.3250 0.3200 1.5550 0.3800 ;
        RECT 5.5000 0.3200 5.6700 0.9000 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0600 0.1800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.2500 1.8400 1.3500 ;
        RECT 1.6150 1.1750 1.8400 1.2500 ;
        RECT 1.6150 0.7500 1.7050 1.1750 ;
        RECT 1.6150 0.6600 2.2050 0.7500 ;
        RECT 2.1150 0.7500 2.2050 1.6500 ;
        RECT 2.1150 1.6500 3.2550 1.7400 ;
    END
    ANTENNAGATEAREA 0.1026 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 1.1650 5.5500 1.4000 ;
        RECT 5.4500 1.0750 5.7100 1.1650 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.3500 4.7500 1.7200 ;
        RECT 4.1350 1.2500 4.7500 1.3500 ;
        RECT 4.1350 1.3500 4.2350 1.7200 ;
        RECT 4.6500 0.9500 4.7500 1.2500 ;
        RECT 4.1400 0.8500 4.7500 0.9500 ;
        RECT 4.1400 0.7050 4.2300 0.8500 ;
        RECT 4.6500 0.7050 4.7500 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 1.6150 2.0100 1.7850 2.0800 ;
        RECT 0.0900 1.6600 0.1800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3500 0.5150 0.4400 1.9300 ;
      RECT 1.3150 1.0500 1.5250 1.1400 ;
      RECT 0.5700 1.5450 0.8650 1.6350 ;
      RECT 0.7750 0.9150 0.8650 1.5450 ;
      RECT 0.7750 0.8250 1.4050 0.9150 ;
      RECT 1.3150 0.9150 1.4050 1.0500 ;
      RECT 1.0900 1.6400 2.0250 1.7300 ;
      RECT 1.9350 0.9300 2.0250 1.6400 ;
      RECT 1.8150 0.8400 2.0250 0.9300 ;
      RECT 1.0900 1.2100 1.1800 1.6400 ;
      RECT 2.3000 1.4600 3.3000 1.5500 ;
      RECT 3.2100 1.1700 3.3000 1.4600 ;
      RECT 2.3000 0.7350 2.3900 1.4600 ;
      RECT 3.2100 1.0800 3.7400 1.1700 ;
      RECT 3.8650 1.0500 4.5150 1.1400 ;
      RECT 3.5600 1.6300 3.9550 1.7200 ;
      RECT 3.8650 1.1400 3.9550 1.6300 ;
      RECT 3.8650 0.8500 3.9550 1.0500 ;
      RECT 2.7650 0.7600 3.9550 0.8500 ;
      RECT 2.7650 0.8500 2.8550 1.3450 ;
      RECT 0.5400 0.4800 5.3200 0.5700 ;
      RECT 5.2300 0.5700 5.3200 1.4700 ;
      RECT 2.5050 0.5700 2.5950 1.3700 ;
      RECT 0.5400 0.5700 0.6300 1.4200 ;
      RECT 5.0400 1.7000 5.8900 1.7900 ;
      RECT 5.8000 0.5250 5.8900 1.7000 ;
      RECT 0.7100 1.8300 5.1400 1.9200 ;
      RECT 5.0400 1.7900 5.1400 1.8300 ;
      RECT 5.0400 1.0050 5.1400 1.7000 ;
      RECT 2.4400 1.9200 2.6100 1.9800 ;
  END
END DFFSQ_X4M_A12TH

MACRO DFFSRPQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8900 ;
        RECT 2.6350 0.3200 2.9250 0.3850 ;
        RECT 5.5300 0.3200 5.6200 0.7700 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 1.1550 5.5500 1.3900 ;
        RECT 5.4500 1.0450 5.7350 1.1550 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 0.9000 2.0600 1.2700 2.0800 ;
        RECT 0.0800 1.5250 0.1700 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8100 5.1500 1.5700 ;
        RECT 4.6900 1.5700 5.1500 1.6600 ;
        RECT 4.6900 0.7200 5.1500 0.8100 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8100 1.0450 4.1400 1.1750 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END R

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0800 3.0700 1.2500 ;
        RECT 2.8500 1.0100 2.9500 1.0800 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0450 0.1600 1.4300 ;
    END
    ANTENNAGATEAREA 0.0192 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6800 0.4300 1.7350 ;
      RECT 0.5550 1.6000 0.7900 1.6900 ;
      RECT 0.7000 1.1900 0.7900 1.6000 ;
      RECT 0.7000 1.1000 1.3450 1.1900 ;
      RECT 1.2550 1.1900 1.3450 1.2850 ;
      RECT 0.7000 0.6800 0.7900 1.1000 ;
      RECT 1.2550 1.2850 1.7800 1.3750 ;
      RECT 1.5450 1.0800 2.1000 1.1700 ;
      RECT 2.0100 0.9300 2.1000 1.0800 ;
      RECT 1.5450 0.7800 1.6350 1.0800 ;
      RECT 2.0100 0.8400 2.2050 0.9300 ;
      RECT 0.9950 1.6000 2.4050 1.6900 ;
      RECT 0.9950 1.2800 1.0850 1.6000 ;
      RECT 2.3150 0.7500 2.4050 1.6000 ;
      RECT 1.8050 0.6600 2.4050 0.7500 ;
      RECT 1.8050 0.7500 1.8950 0.9900 ;
      RECT 3.3700 0.6600 4.3400 0.7500 ;
      RECT 4.2500 0.7500 4.3400 1.3750 ;
      RECT 2.5400 1.6400 3.4600 1.7300 ;
      RECT 3.3700 0.7500 3.4600 1.6400 ;
      RECT 2.5400 0.8750 2.6300 1.6400 ;
      RECT 2.5400 0.7850 2.7300 0.8750 ;
      RECT 4.4750 1.2000 4.9300 1.2900 ;
      RECT 3.7500 1.6400 4.5650 1.7300 ;
      RECT 3.7500 1.3500 3.8400 1.6400 ;
      RECT 4.4750 1.2900 4.5650 1.6400 ;
      RECT 4.4750 0.6600 4.5650 1.2000 ;
      RECT 0.5200 0.4800 5.3300 0.5700 ;
      RECT 5.2400 0.5700 5.3300 1.7200 ;
      RECT 3.1700 0.5700 3.2600 1.5500 ;
      RECT 0.5200 0.5700 0.6100 1.4900 ;
      RECT 0.6600 1.8300 5.9150 1.9200 ;
      RECT 5.8250 1.7150 5.9150 1.8300 ;
      RECT 5.8250 1.6550 5.9200 1.7150 ;
      RECT 5.8300 0.5600 5.9200 1.6550 ;
      RECT 3.5600 0.8850 3.6500 1.8300 ;
  END
END DFFSRPQ_X0P5M_A12TH

MACRO DFFSRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7950 ;
        RECT 5.4700 0.3200 5.6400 0.8150 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6400 0.9550 5.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.9500 4.9500 1.2500 ;
        RECT 4.8500 1.2500 5.0850 1.3500 ;
        RECT 4.8500 0.8500 5.0850 0.9500 ;
        RECT 4.9950 1.3500 5.0850 1.7100 ;
        RECT 4.9950 0.7050 5.0850 0.8500 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0000 1.0100 4.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0588 ;
  END R

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9800 0.1600 1.4050 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0400 0.9600 3.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END SN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 0.0800 1.5250 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.7050 0.4300 1.7650 ;
      RECT 0.5800 1.5900 0.7900 1.6800 ;
      RECT 0.7000 1.1450 0.7900 1.5900 ;
      RECT 0.7000 1.0550 1.3650 1.1450 ;
      RECT 1.2750 1.1450 1.3650 1.2300 ;
      RECT 0.7000 0.6800 0.7900 1.0550 ;
      RECT 1.2750 1.2300 1.7600 1.3200 ;
      RECT 1.6700 1.3200 1.7600 1.4600 ;
      RECT 1.5700 1.0050 2.1200 1.0950 ;
      RECT 2.0300 0.9300 2.1200 1.0050 ;
      RECT 1.5700 0.7800 1.6600 1.0050 ;
      RECT 2.0300 0.8400 2.2400 0.9300 ;
      RECT 0.9950 1.5700 2.4500 1.6600 ;
      RECT 0.9950 1.2550 1.0850 1.5700 ;
      RECT 2.3600 0.7500 2.4500 1.5700 ;
      RECT 1.8300 0.6600 2.4500 0.7500 ;
      RECT 1.8300 0.7500 1.9200 0.9150 ;
      RECT 3.4300 0.6700 4.4250 0.7600 ;
      RECT 4.3350 0.7600 4.4250 1.3450 ;
      RECT 2.6650 1.6450 3.5200 1.7350 ;
      RECT 3.4300 0.7600 3.5200 1.6450 ;
      RECT 2.6650 1.5850 2.7550 1.6450 ;
      RECT 2.5400 1.4950 2.7550 1.5850 ;
      RECT 2.6650 0.8950 2.7550 1.4950 ;
      RECT 2.5600 0.8050 2.7550 0.8950 ;
      RECT 3.8200 1.6400 4.6200 1.7300 ;
      RECT 4.5300 1.1550 4.6200 1.6400 ;
      RECT 4.5300 1.0650 4.7600 1.1550 ;
      RECT 4.5300 0.6800 4.6200 1.0650 ;
      RECT 3.8200 1.3500 3.9100 1.6400 ;
      RECT 0.5200 0.4800 5.3150 0.5700 ;
      RECT 5.2250 0.5700 5.3150 1.5700 ;
      RECT 3.2400 0.5700 3.3300 1.5350 ;
      RECT 0.5200 0.5700 0.6100 1.4750 ;
      RECT 5.5300 1.4800 5.9450 1.5700 ;
      RECT 5.8550 0.8300 5.9450 1.4800 ;
      RECT 5.7550 0.7400 5.9450 0.8300 ;
      RECT 0.7000 1.8300 5.6200 1.9200 ;
      RECT 5.5300 1.5700 5.6200 1.8300 ;
      RECT 3.6300 0.8500 3.7200 1.8300 ;
  END
END DFFSRPQ_X1M_A12TH

MACRO DFFSRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8400 ;
        RECT 5.6650 0.3200 5.8350 0.7600 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.1600 5.7500 1.3900 ;
        RECT 5.6500 1.0500 5.9100 1.1600 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 4.2050 2.0350 4.3450 2.0800 ;
        RECT 5.6700 1.8850 5.8400 2.0800 ;
        RECT 0.0800 1.5950 0.1700 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8450 5.1500 1.2500 ;
        RECT 4.9550 1.2500 5.1500 1.3500 ;
        RECT 4.8950 0.7550 5.1500 0.8450 ;
        RECT 4.9550 1.3500 5.0450 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1800 4.1500 1.3900 ;
        RECT 3.8700 1.0900 4.1500 1.1800 ;
    END
    ANTENNAGATEAREA 0.0714 ;
  END R

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.2000 2.9500 1.3900 ;
        RECT 2.8500 1.1000 3.1350 1.2000 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.4650 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6300 0.4300 1.7650 ;
      RECT 0.5450 1.5900 0.7900 1.6800 ;
      RECT 0.7000 1.1750 0.7900 1.5900 ;
      RECT 0.7000 1.0850 1.7600 1.1750 ;
      RECT 1.6700 1.1750 1.7600 1.2750 ;
      RECT 0.7000 0.6800 0.7900 1.0850 ;
      RECT 1.5100 0.6750 2.2400 0.7650 ;
      RECT 1.0550 1.5700 2.4450 1.6600 ;
      RECT 1.0550 1.2650 1.1450 1.5700 ;
      RECT 2.3550 0.9550 2.4450 1.5700 ;
      RECT 1.7700 0.8650 2.4450 0.9550 ;
      RECT 2.3550 0.7550 2.4450 0.8650 ;
      RECT 3.4050 0.6600 4.4000 0.7500 ;
      RECT 4.3100 0.7500 4.4000 1.4200 ;
      RECT 2.5350 1.6450 3.4950 1.7350 ;
      RECT 3.4050 0.7500 3.4950 1.6450 ;
      RECT 2.5350 0.8950 2.6250 1.6450 ;
      RECT 2.5350 0.8050 2.7800 0.8950 ;
      RECT 3.7950 1.6400 4.5800 1.7300 ;
      RECT 4.4900 1.1700 4.5800 1.6400 ;
      RECT 4.4900 1.0800 4.7450 1.1700 ;
      RECT 4.4900 0.7050 4.5800 1.0800 ;
      RECT 3.7950 1.3500 3.8850 1.6400 ;
      RECT 0.5200 0.4800 5.5100 0.5700 ;
      RECT 5.4200 0.5700 5.5100 1.5600 ;
      RECT 3.2250 0.5700 3.3150 1.5350 ;
      RECT 0.5200 0.5700 0.6100 1.4750 ;
      RECT 5.4450 1.6550 6.0900 1.7450 ;
      RECT 6.0000 0.6050 6.0900 1.6550 ;
      RECT 0.7100 1.8300 5.5350 1.9200 ;
      RECT 5.4450 1.7450 5.5350 1.8300 ;
      RECT 3.6050 0.8650 3.6950 1.8300 ;
  END
END DFFSRPQ_X2M_A12TH

MACRO DFFSRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8400 ;
        RECT 2.7500 0.3200 2.9450 0.3700 ;
        RECT 4.2200 0.3200 4.3900 0.3900 ;
        RECT 6.0750 0.3200 6.2450 0.6900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2450 0.8950 6.3650 1.3050 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 1.2000 2.0100 1.3700 2.0800 ;
        RECT 1.9450 2.0100 2.1150 2.0800 ;
        RECT 0.0800 1.6950 0.1700 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0850 0.8500 5.6950 0.9500 ;
        RECT 5.4500 0.9500 5.5500 1.2500 ;
        RECT 5.0850 0.6850 5.1750 0.8500 ;
        RECT 5.6050 0.6850 5.6950 0.8500 ;
        RECT 5.0850 1.2500 5.6950 1.3500 ;
        RECT 5.0850 1.3500 5.1750 1.7200 ;
        RECT 5.6050 1.3500 5.6950 1.7200 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0500 1.9700 1.4350 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END R

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 1.0050 3.9500 1.2200 ;
        RECT 3.8500 0.9050 4.1200 1.0050 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0450 0.1800 1.4150 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 0.5000 0.4300 1.9850 ;
      RECT 0.5450 1.5900 0.7900 1.6800 ;
      RECT 0.7000 1.1500 0.7900 1.5900 ;
      RECT 0.7000 1.0600 1.6950 1.1500 ;
      RECT 1.6050 1.1500 1.6950 1.2950 ;
      RECT 0.7000 0.6800 0.7900 1.0600 ;
      RECT 1.4550 0.6700 2.1850 0.7600 ;
      RECT 0.9950 1.6400 2.4150 1.7300 ;
      RECT 2.3250 0.9400 2.4150 1.6400 ;
      RECT 1.7150 0.8500 2.4150 0.9400 ;
      RECT 0.9950 1.2400 1.0850 1.6400 ;
      RECT 3.3800 0.6700 4.4300 0.7600 ;
      RECT 4.3400 0.7600 4.4300 1.1250 ;
      RECT 2.5450 1.6450 3.4700 1.7350 ;
      RECT 2.5450 0.7750 2.6350 1.6450 ;
      RECT 3.3800 0.7600 3.4700 1.6450 ;
      RECT 4.5200 1.0650 5.3400 1.1550 ;
      RECT 3.7400 1.6500 4.6100 1.7400 ;
      RECT 4.5200 1.1550 4.6100 1.6500 ;
      RECT 4.5200 0.7600 4.6100 1.0650 ;
      RECT 4.5200 0.6700 4.6900 0.7600 ;
      RECT 3.7400 1.3700 3.8300 1.6500 ;
      RECT 0.5200 0.4800 5.9450 0.5700 ;
      RECT 5.8550 0.5700 5.9450 1.6100 ;
      RECT 3.2000 0.5700 3.2900 1.5350 ;
      RECT 2.4300 0.4100 2.6000 0.4800 ;
      RECT 0.5200 0.5700 0.6100 1.4750 ;
      RECT 6.0350 1.5450 6.5550 1.6350 ;
      RECT 6.4650 0.6650 6.5550 1.5450 ;
      RECT 6.3450 0.5750 6.5550 0.6650 ;
      RECT 0.7000 1.8300 6.1250 1.9200 ;
      RECT 6.0350 1.6350 6.1250 1.8300 ;
      RECT 6.0350 0.9800 6.1250 1.5450 ;
      RECT 2.4300 1.9200 2.6000 1.9800 ;
      RECT 3.5600 0.8850 3.6500 1.8300 ;
  END
END DFFSRPQ_X3M_A12TH

MACRO DFFSRPQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6800 ;
        RECT 6.2950 0.3200 6.4650 0.5350 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4450 0.9150 6.5500 1.3350 ;
    END
    ANTENNAGATEAREA 0.033 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 0.0950 1.7600 0.1850 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0450 0.8500 5.7500 0.9500 ;
        RECT 5.6500 0.9500 5.7500 1.2500 ;
        RECT 5.0450 0.7050 5.1350 0.8500 ;
        RECT 5.5650 0.7050 5.6550 0.8500 ;
        RECT 5.0450 1.2500 5.7500 1.3500 ;
        RECT 5.0450 1.3500 5.1350 1.7150 ;
        RECT 5.5650 1.3500 5.6550 1.7150 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.8800 4.1500 1.1100 ;
        RECT 3.9250 1.1100 4.1500 1.2100 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END R

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 1.0500 3.1700 1.4500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END SN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0450 0.1600 1.4300 ;
    END
    ANTENNAGATEAREA 0.0768 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3550 0.4300 0.4450 1.9500 ;
      RECT 0.5550 1.5650 0.8250 1.6550 ;
      RECT 0.7350 0.9600 0.8250 1.5650 ;
      RECT 0.7350 0.8700 1.6300 0.9600 ;
      RECT 1.5400 0.9600 1.6300 1.1400 ;
      RECT 0.7350 0.6800 0.8250 0.8700 ;
      RECT 1.5400 1.1400 1.8050 1.2300 ;
      RECT 1.4900 0.6700 2.2200 0.7600 ;
      RECT 1.0950 1.6400 2.0100 1.7300 ;
      RECT 1.0950 1.0550 1.1850 1.6400 ;
      RECT 1.9200 0.9400 2.0100 1.6400 ;
      RECT 1.7500 0.8500 2.4950 0.9400 ;
      RECT 2.4050 0.9400 2.4950 1.5200 ;
      RECT 2.3600 1.5200 2.4950 1.6900 ;
      RECT 3.4550 0.6700 4.3550 0.7600 ;
      RECT 4.2650 0.7600 4.3550 1.1950 ;
      RECT 4.2650 1.1950 4.7600 1.2850 ;
      RECT 2.6200 1.6450 3.5450 1.7350 ;
      RECT 3.4550 0.7600 3.5450 1.6450 ;
      RECT 2.6200 0.7450 2.7100 1.6450 ;
      RECT 4.8500 1.0650 5.4400 1.1550 ;
      RECT 3.8400 1.6400 4.9400 1.7300 ;
      RECT 4.8500 1.1550 4.9400 1.6400 ;
      RECT 4.8500 0.7700 4.9400 1.0650 ;
      RECT 4.4650 0.6800 4.9400 0.7700 ;
      RECT 3.8400 1.3500 3.9300 1.6400 ;
      RECT 0.5550 0.4800 6.1650 0.5700 ;
      RECT 6.0750 0.5700 6.1650 1.5200 ;
      RECT 3.2600 0.5700 3.3500 1.5300 ;
      RECT 0.5550 0.5700 0.6450 1.4550 ;
      RECT 2.8000 0.5700 2.8900 1.1600 ;
      RECT 0.7600 1.8300 6.4900 1.9200 ;
      RECT 6.4000 1.5900 6.4900 1.8300 ;
      RECT 6.4000 1.5000 6.7350 1.5900 ;
      RECT 6.6450 0.7250 6.7350 1.5000 ;
      RECT 6.2550 0.6350 6.7350 0.7250 ;
      RECT 6.6300 0.4450 6.7350 0.6350 ;
      RECT 6.2550 0.7250 6.3450 0.9350 ;
      RECT 3.6550 0.8700 3.7450 1.8300 ;
      RECT 2.1750 1.2200 2.2650 1.8300 ;
  END
END DFFSRPQ_X4M_A12TH

MACRO DFFYQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8050 ;
        RECT 1.2350 0.3200 1.4050 0.4800 ;
        RECT 2.5350 0.3200 2.6250 0.3900 ;
        RECT 3.3350 0.3200 3.5050 0.3750 ;
        RECT 3.7650 0.3200 3.8650 0.5500 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.8900 3.9500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9500 3.1500 1.3100 ;
        RECT 2.9450 1.3100 3.1500 1.4100 ;
        RECT 3.0500 0.8500 3.1950 0.9500 ;
        RECT 2.9450 1.4100 3.0450 1.7200 ;
        RECT 3.0950 0.7450 3.1950 0.8500 ;
    END
    ANTENNADIFFAREA 0.26455 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 2.2900 2.0300 2.4600 2.0800 ;
        RECT 1.1300 2.0100 1.3000 2.0800 ;
        RECT 0.0800 1.7750 0.1700 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2200 0.1700 1.4200 ;
        RECT 0.0500 1.0500 0.2300 1.2200 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.3400 0.5950 0.4300 1.7550 ;
      RECT 0.5750 1.6100 0.7950 1.7000 ;
      RECT 0.7050 1.4300 0.7950 1.6100 ;
      RECT 0.7050 1.3400 1.4550 1.4300 ;
      RECT 0.7050 0.6800 0.7950 1.3400 ;
      RECT 1.5450 1.2200 1.6350 1.7200 ;
      RECT 1.0050 1.1300 1.6350 1.2200 ;
      RECT 1.5450 0.8450 1.6350 1.1300 ;
      RECT 1.5450 0.7550 1.7500 0.8450 ;
      RECT 1.7450 1.5600 1.9500 1.6500 ;
      RECT 1.8600 0.7850 1.9500 1.5600 ;
      RECT 1.8600 0.6950 2.4800 0.7850 ;
      RECT 2.3900 0.7850 2.4800 0.8850 ;
      RECT 2.3900 0.8850 2.6950 0.9950 ;
      RECT 2.8150 0.6600 2.9850 0.7500 ;
      RECT 2.2200 1.6200 2.8050 1.7100 ;
      RECT 2.2200 1.2800 2.3100 1.6200 ;
      RECT 2.7150 1.2150 2.8050 1.6200 ;
      RECT 2.7150 1.0850 2.9050 1.2150 ;
      RECT 2.8150 0.7500 2.9050 1.0850 ;
      RECT 3.3050 1.4950 3.6900 1.5850 ;
      RECT 3.3050 0.9000 3.3950 1.4950 ;
      RECT 3.3050 0.8100 3.7500 0.9000 ;
      RECT 3.6600 0.7050 3.7500 0.8100 ;
      RECT 3.3050 0.5700 3.3950 0.8100 ;
      RECT 1.6450 0.4800 3.3950 0.5700 ;
      RECT 0.9050 0.5700 1.7350 0.6600 ;
      RECT 1.7850 0.4100 1.9550 0.4800 ;
      RECT 0.9050 0.6600 0.9950 1.0300 ;
      RECT 0.5250 0.4800 0.9950 0.5700 ;
      RECT 0.5250 0.5700 0.6150 1.5000 ;
      RECT 3.4650 1.7000 4.1400 1.7900 ;
      RECT 4.0300 1.5800 4.1400 1.7000 ;
      RECT 4.0500 0.6000 4.1400 1.5800 ;
      RECT 3.9950 0.4300 4.1400 0.6000 ;
      RECT 0.7100 1.9200 0.8800 1.9900 ;
      RECT 0.7100 1.8300 3.5550 1.9200 ;
      RECT 3.4650 1.7900 3.5550 1.8300 ;
      RECT 1.5800 1.9200 1.7500 1.9900 ;
      RECT 2.0400 1.1500 2.1300 1.8300 ;
      RECT 2.0400 1.0600 2.2700 1.1500 ;
  END
END DFFYQ_X1M_A12TH

MACRO DFFYQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.4250 0.3200 0.5150 0.4500 ;
        RECT 0.9050 0.3200 1.0750 0.5250 ;
        RECT 2.3300 0.3200 2.4200 0.5650 ;
        RECT 3.6100 0.3200 3.7000 0.8900 ;
        RECT 4.4300 0.3200 4.5200 0.5000 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3900 1.2100 4.5500 1.4250 ;
        RECT 4.3900 1.0900 4.4800 1.2100 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9150 0.9500 1.5250 ;
        RECT 0.6800 1.5250 0.9500 1.6250 ;
        RECT 0.6250 0.8150 0.9500 0.9150 ;
        RECT 0.6800 1.6250 0.7800 1.9350 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.1800 3.5500 1.6000 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 4.4300 1.9000 4.5200 2.0800 ;
        RECT 0.9450 1.7700 1.0350 2.0800 ;
        RECT 0.4100 1.6900 0.5000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.3450 0.7200 1.4350 ;
      RECT 0.6300 1.0250 0.7200 1.3450 ;
      RECT 0.0800 1.4350 0.1700 1.7550 ;
      RECT 0.0800 0.5250 0.1700 1.3450 ;
      RECT 1.5100 1.6750 1.6000 1.8050 ;
      RECT 1.1500 1.5850 1.6000 1.6750 ;
      RECT 1.1500 0.7050 1.2400 1.5850 ;
      RECT 0.2600 0.6150 1.6200 0.7050 ;
      RECT 1.5300 0.4950 1.6200 0.6150 ;
      RECT 0.2600 0.7050 0.3550 1.2150 ;
      RECT 1.8900 1.6000 2.5450 1.6900 ;
      RECT 2.4550 1.3250 2.5450 1.6000 ;
      RECT 1.8900 0.8050 1.9800 1.6000 ;
      RECT 1.8900 0.7150 2.0600 0.8050 ;
      RECT 2.7100 1.6050 2.9400 1.6950 ;
      RECT 2.7100 1.2350 2.8000 1.6050 ;
      RECT 2.1050 1.1450 2.8000 1.2350 ;
      RECT 2.1050 1.0250 2.1950 1.1450 ;
      RECT 2.7100 0.7750 2.8000 1.1450 ;
      RECT 2.7100 0.6850 2.9800 0.7750 ;
      RECT 3.2500 0.6800 3.3400 1.7400 ;
      RECT 1.7100 1.8300 4.0300 1.9200 ;
      RECT 3.9400 1.7650 4.0300 1.8300 ;
      RECT 3.9400 1.5550 4.0800 1.7650 ;
      RECT 3.9900 0.7750 4.0800 1.5550 ;
      RECT 3.0500 1.5150 3.1400 1.8300 ;
      RECT 1.7100 1.4950 1.8000 1.8300 ;
      RECT 2.8900 1.4250 3.1400 1.5150 ;
      RECT 1.3800 1.4050 1.8000 1.4950 ;
      RECT 2.8900 0.8850 2.9800 1.4250 ;
      RECT 1.7100 1.0850 1.8000 1.4050 ;
      RECT 1.5850 0.9950 1.8000 1.0850 ;
      RECT 3.7850 1.0900 3.8800 1.2000 ;
      RECT 3.4300 1.0000 3.8800 1.0900 ;
      RECT 3.7900 0.6650 3.8800 1.0000 ;
      RECT 3.7900 0.5750 4.2600 0.6650 ;
      RECT 4.1700 0.6650 4.2600 1.9650 ;
      RECT 4.1700 0.4100 4.2600 0.5750 ;
      RECT 2.1500 0.6050 2.2400 0.7050 ;
      RECT 1.7100 0.5150 2.2400 0.6050 ;
      RECT 1.7100 0.6050 1.8000 0.8150 ;
      RECT 1.3850 0.8150 1.8000 0.9050 ;
      RECT 1.3850 0.9050 1.4750 1.2750 ;
      RECT 3.4300 0.5700 3.5200 1.0000 ;
      RECT 2.5300 0.4800 3.5200 0.5700 ;
      RECT 2.5300 0.5700 2.6200 0.7050 ;
      RECT 3.0700 0.5700 3.1600 1.3150 ;
      RECT 2.1500 0.7050 2.6200 0.7950 ;
  END
END DFFYQ_X2M_A12TH

MACRO DFFYQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6400 ;
        RECT 0.8600 0.3200 0.9700 0.4400 ;
        RECT 4.1100 0.3200 4.3150 0.3800 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8100 1.0500 0.9900 ;
        RECT 0.9600 0.9900 1.0500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0432 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0800 1.2100 4.3500 1.4200 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4500 0.6900 1.5500 ;
        RECT 0.0500 1.5500 0.1800 1.8800 ;
        RECT 0.6000 1.5500 0.6900 1.8850 ;
        RECT 0.0500 0.9200 0.1500 1.4500 ;
        RECT 0.0500 0.8200 0.6950 0.9200 ;
        RECT 0.0500 0.4900 0.1750 0.8200 ;
        RECT 0.5950 0.4900 0.6950 0.8200 ;
    END
    ANTENNADIFFAREA 0.593125 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 4.0350 2.0150 4.2450 2.0800 ;
        RECT 0.8600 1.8200 0.9600 2.0800 ;
        RECT 0.3350 1.8000 0.4350 2.0800 ;
        RECT 1.7150 1.7200 1.8050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.3400 0.8800 1.9450 0.9700 ;
      RECT 0.7800 1.6400 1.5000 1.7300 ;
      RECT 1.3400 1.3200 1.5000 1.6400 ;
      RECT 1.3400 0.9700 1.4300 1.3200 ;
      RECT 1.3400 0.6600 1.4300 0.8800 ;
      RECT 0.7800 1.1800 0.8700 1.6400 ;
      RECT 0.3750 1.0900 0.8700 1.1800 ;
      RECT 1.9700 1.8750 2.3850 1.9650 ;
      RECT 1.9700 1.5650 2.0600 1.8750 ;
      RECT 1.8000 1.4750 2.0600 1.5650 ;
      RECT 1.8000 1.1850 1.8900 1.4750 ;
      RECT 1.5200 1.1500 1.8900 1.1850 ;
      RECT 1.5200 1.0950 2.2400 1.1500 ;
      RECT 1.8000 1.0600 2.2400 1.0950 ;
      RECT 2.1500 0.7700 2.2400 1.0600 ;
      RECT 2.1500 0.6800 2.3450 0.7700 ;
      RECT 2.6000 1.4950 2.7900 1.5850 ;
      RECT 2.7000 1.3450 2.7900 1.4950 ;
      RECT 2.7000 1.2550 3.0900 1.3450 ;
      RECT 3.0000 1.1550 3.0900 1.2550 ;
      RECT 2.7000 0.7700 2.7900 1.2550 ;
      RECT 2.6150 0.6800 2.7900 0.7700 ;
      RECT 3.4500 1.4250 3.5500 1.7200 ;
      RECT 3.2000 1.3350 3.5500 1.4250 ;
      RECT 3.2000 0.8900 3.2900 1.3350 ;
      RECT 2.9000 0.8000 3.5900 0.8900 ;
      RECT 2.9000 0.8900 2.9900 1.0550 ;
      RECT 3.5000 0.6600 3.5900 0.8000 ;
      RECT 3.8350 1.5700 3.9900 1.7400 ;
      RECT 3.9000 0.6600 3.9900 1.5700 ;
      RECT 1.1400 0.4800 4.2000 0.5700 ;
      RECT 4.1100 0.5700 4.2000 0.8600 ;
      RECT 4.1100 0.8600 4.3500 0.9500 ;
      RECT 4.2600 0.9500 4.3500 1.0700 ;
      RECT 2.0000 1.2400 2.5650 1.3300 ;
      RECT 2.4350 1.1600 2.5650 1.2400 ;
      RECT 2.4350 0.5700 2.5250 1.1600 ;
      RECT 1.1400 0.5700 1.2300 1.5100 ;
      RECT 3.7000 0.5700 3.7900 1.0650 ;
      RECT 1.1400 0.4100 1.3150 0.4800 ;
      RECT 3.1050 1.8300 4.5300 1.9200 ;
      RECT 4.4400 0.6350 4.5300 1.8300 ;
      RECT 4.4300 0.4100 4.5300 0.6350 ;
      RECT 3.1050 1.7750 3.1950 1.8300 ;
      RECT 3.6400 1.2450 3.7350 1.8300 ;
      RECT 2.2300 1.6850 3.1950 1.7750 ;
      RECT 3.5000 1.1550 3.7350 1.2450 ;
      RECT 2.2300 1.6050 2.3200 1.6850 ;
      RECT 3.5000 1.0800 3.5900 1.1550 ;
      RECT 2.1500 1.5150 2.3200 1.6050 ;
      RECT 3.4000 0.9800 3.5900 1.0800 ;
  END
END DFFYQ_X3M_A12TH

MACRO DFFYQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.4050 0.3200 0.4950 0.4700 ;
        RECT 0.9250 0.3200 1.0150 0.4700 ;
        RECT 1.4450 0.3200 1.5350 0.4700 ;
        RECT 1.9700 0.3200 2.0600 0.4700 ;
        RECT 3.3350 0.3200 3.5450 0.4200 ;
        RECT 4.7300 0.3200 4.8200 0.3900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 0.9200 0.3500 1.2900 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6000 1.4500 1.2200 1.5500 ;
        RECT 0.6000 1.5500 0.7000 1.8550 ;
        RECT 1.1200 1.5500 1.2200 1.8550 ;
        RECT 0.6500 0.9500 0.7550 1.4500 ;
        RECT 0.6500 0.8500 1.2800 0.9500 ;
        RECT 0.6500 0.7700 0.7600 0.8500 ;
        RECT 1.1800 0.7700 1.2800 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.1000 4.7500 1.5200 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 4.7000 2.0100 4.8950 2.0800 ;
        RECT 3.5550 1.8300 3.6450 2.0800 ;
        RECT 0.8650 1.7700 0.9550 2.0800 ;
        RECT 1.3850 1.7700 1.4750 2.0800 ;
        RECT 1.6350 1.7500 1.7250 2.0800 ;
        RECT 2.2150 1.7500 2.3050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.9200 1.0500 2.2400 1.0650 ;
      RECT 2.1500 1.0650 2.2400 1.1850 ;
      RECT 1.4550 0.9750 2.2400 1.0500 ;
      RECT 1.4550 1.1400 1.5450 1.5150 ;
      RECT 0.9200 1.0650 1.5450 1.1400 ;
      RECT 1.8950 1.6050 1.9850 1.9450 ;
      RECT 1.4550 1.5150 1.9850 1.6050 ;
      RECT 1.7100 0.7700 1.8000 0.9750 ;
      RECT 2.7850 1.6000 2.8750 1.9650 ;
      RECT 2.3400 1.5100 2.8750 1.6000 ;
      RECT 2.3400 1.4050 2.4300 1.5100 ;
      RECT 1.7300 1.3150 2.4300 1.4050 ;
      RECT 2.3400 0.8600 2.4300 1.3150 ;
      RECT 2.3400 0.7700 2.7300 0.8600 ;
      RECT 2.5600 0.7100 2.7300 0.7700 ;
      RECT 3.1650 0.9700 3.2550 1.6600 ;
      RECT 3.1650 0.8700 3.6000 0.9700 ;
      RECT 3.1650 0.8000 3.2550 0.8700 ;
      RECT 3.0000 0.7100 3.2550 0.8000 ;
      RECT 4.1100 1.5350 4.2000 1.7200 ;
      RECT 3.6900 1.4450 4.2000 1.5350 ;
      RECT 3.6900 1.1950 3.7800 1.4450 ;
      RECT 3.3450 1.1050 3.7800 1.1950 ;
      RECT 3.6900 0.8000 3.7800 1.1050 ;
      RECT 3.6900 0.7100 4.1600 0.8000 ;
      RECT 3.9700 0.6600 4.1600 0.7100 ;
      RECT 4.4700 0.6600 4.5600 1.7200 ;
      RECT 2.2700 0.5100 4.7600 0.5700 ;
      RECT 4.6700 0.5700 4.7600 0.9000 ;
      RECT 3.7000 0.4800 4.7600 0.5100 ;
      RECT 4.6700 0.9000 4.9300 0.9900 ;
      RECT 4.8400 0.9900 4.9300 1.1700 ;
      RECT 0.4500 0.6000 2.3600 0.6800 ;
      RECT 0.4500 0.5900 3.7900 0.6000 ;
      RECT 2.8200 0.6000 2.9100 1.0500 ;
      RECT 2.2700 0.5700 3.7900 0.5900 ;
      RECT 2.5200 1.0500 3.0550 1.1400 ;
      RECT 2.9650 1.1400 3.0550 1.2200 ;
      RECT 2.5200 0.9700 2.6100 1.0500 ;
      RECT 4.2700 0.5700 4.3600 1.1350 ;
      RECT 0.0800 1.4700 0.1700 1.7500 ;
      RECT 0.0500 1.3800 0.1700 1.4700 ;
      RECT 0.0500 0.8300 0.1400 1.3800 ;
      RECT 0.0800 0.4600 0.1700 0.7400 ;
      RECT 0.0500 0.7400 0.5400 0.8300 ;
      RECT 0.4500 0.6800 0.5400 0.7400 ;
      RECT 3.8500 1.8300 5.1200 1.9200 ;
      RECT 5.0300 0.4900 5.1200 1.8300 ;
      RECT 3.8500 1.7350 3.9400 1.8300 ;
      RECT 4.2900 1.3350 4.3800 1.8300 ;
      RECT 3.3550 1.6450 3.9400 1.7350 ;
      RECT 4.0900 1.2450 4.3800 1.3350 ;
      RECT 4.0900 0.9800 4.1800 1.2450 ;
      RECT 3.8900 0.8900 4.1800 0.9800 ;
      RECT 3.3550 1.7350 3.4450 1.7700 ;
      RECT 2.9650 1.7700 3.4450 1.8600 ;
      RECT 2.9650 1.4100 3.0550 1.7700 ;
      RECT 2.6250 1.3200 3.0550 1.4100 ;
  END
END DFFYQ_X4M_A12TH

MACRO DLY2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3850 0.3200 0.4750 0.6100 ;
        RECT 0.7250 0.3200 0.8150 0.8100 ;
        RECT 0.9800 0.3200 1.0800 0.4900 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9850 1.8850 1.0750 2.0800 ;
        RECT 0.3850 1.6700 0.4750 2.0800 ;
        RECT 0.7250 1.3200 0.8150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8450 1.1500 1.2900 ;
        RECT 0.9850 1.2900 1.1500 1.7000 ;
        RECT 0.9250 0.7550 1.1500 0.8450 ;
    END
    ANTENNADIFFAREA 0.16605 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0100 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0432 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.1250 1.3200 0.2150 1.8800 ;
      RECT 0.1250 0.4200 0.2150 0.9000 ;
      RECT 0.4950 1.0750 0.9000 1.1650 ;
      RECT 0.3250 1.3800 0.5850 1.4700 ;
      RECT 0.4950 1.1650 0.5850 1.3800 ;
      RECT 0.4950 0.8400 0.5850 1.0750 ;
      RECT 0.3250 0.7500 0.5850 0.8400 ;
  END
END DLY2_X0P5M_A12TH

MACRO DLY2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.7500 1.7700 0.8500 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.7500 0.3200 0.8500 0.6500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9150 1.1500 1.2900 ;
        RECT 1.0300 1.2900 1.1500 1.7100 ;
        RECT 1.0250 0.4750 1.1500 0.9150 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.5500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0564 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0700 1.5750 0.2400 1.9900 ;
      RECT 0.0700 0.4100 0.2400 0.7900 ;
      RECT 0.4050 1.5150 0.7850 1.6050 ;
      RECT 0.6950 0.8550 0.7850 1.5150 ;
      RECT 0.4050 0.7650 0.7850 0.8550 ;
      RECT 0.4050 1.6050 0.4950 1.7750 ;
      RECT 0.4050 0.6400 0.4950 0.7650 ;
  END
END DLY2_X1M_A12TH

MACRO DLY2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.6250 1.7600 0.7250 2.0800 ;
        RECT 0.8950 1.7600 0.9950 2.0800 ;
        RECT 1.4150 1.7600 1.5150 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.6250 0.3200 0.7250 0.6500 ;
        RECT 0.8950 0.3200 0.9950 0.6500 ;
        RECT 1.4150 0.3200 1.5150 0.6500 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.2500 ;
        RECT 1.1550 1.2500 1.5500 1.3500 ;
        RECT 1.1550 0.8500 1.5500 0.9500 ;
        RECT 1.1550 1.3500 1.2550 1.7100 ;
        RECT 1.1550 0.4750 1.2550 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.5500 1.1900 ;
    END
    ANTENNAGATEAREA 0.1584 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0500 1.2550 1.1500 ;
      RECT 0.0850 1.6050 0.1850 1.9400 ;
      RECT 0.0500 0.4100 0.2200 0.7650 ;
      RECT 0.0850 1.5050 0.7900 1.6050 ;
      RECT 0.7000 1.1500 0.7900 1.5050 ;
      RECT 0.7000 0.8650 0.7900 1.0500 ;
      RECT 0.0500 0.7650 0.7900 0.8650 ;
  END
END DLY2_X2M_A12TH

MACRO DLY2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.0750 1.7600 0.1750 2.0800 ;
        RECT 1.0550 1.7600 1.1550 2.0800 ;
        RECT 1.3250 1.7600 1.4250 2.0800 ;
        RECT 1.5850 1.7600 1.6850 2.0800 ;
        RECT 2.1050 1.7600 2.2050 2.0800 ;
        RECT 2.6250 1.7600 2.7250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.0500 1.0000 1.1500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9500 2.5500 1.2500 ;
        RECT 1.8450 1.2500 2.5500 1.3500 ;
        RECT 1.8450 0.8500 2.5500 0.9500 ;
        RECT 1.8450 1.3500 1.9450 1.7100 ;
        RECT 2.3650 1.3500 2.4650 1.7100 ;
        RECT 1.8450 0.4750 1.9450 0.8500 ;
        RECT 2.3650 0.4750 2.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6400 ;
        RECT 1.0550 0.3200 1.1550 0.6500 ;
        RECT 1.3250 0.3200 1.4250 0.6500 ;
        RECT 1.5850 0.3200 1.6850 0.6500 ;
        RECT 2.1050 0.3200 2.2050 0.6500 ;
        RECT 2.6250 0.3200 2.7250 0.6500 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.1300 1.0500 2.3400 1.1500 ;
      RECT 0.5650 1.3500 0.6650 1.7400 ;
      RECT 0.5650 0.4100 0.6650 0.7650 ;
      RECT 0.5650 1.2500 1.2200 1.3500 ;
      RECT 1.1300 1.1500 1.2200 1.2500 ;
      RECT 1.1300 0.8650 1.2200 1.0500 ;
      RECT 0.5650 0.7650 1.2200 0.8650 ;
  END
END DLY2_X4M_A12TH

MACRO DLY4_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3600 0.3200 0.4500 0.6200 ;
        RECT 0.9150 0.3200 1.0050 0.6000 ;
        RECT 1.4650 0.3200 1.5550 0.6000 ;
        RECT 1.7550 0.3200 1.8450 0.9950 ;
        RECT 2.0150 0.3200 2.1050 0.4900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0100 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0432 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0100 0.7150 2.1500 1.5500 ;
    END
    ANTENNADIFFAREA 0.14175 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 2.0150 1.8850 2.1050 2.0800 ;
        RECT 0.9150 1.6700 1.0050 2.0800 ;
        RECT 1.4650 1.6650 1.5550 2.0800 ;
        RECT 0.3600 1.6600 0.4500 2.0800 ;
        RECT 1.7550 1.3300 1.8450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1000 1.3150 0.1900 1.8700 ;
      RECT 0.1000 0.4200 0.1900 0.9000 ;
      RECT 0.6550 1.3100 0.7450 1.8700 ;
      RECT 0.6550 0.4200 0.7450 0.9000 ;
      RECT 0.3000 1.3750 0.5300 1.4650 ;
      RECT 0.4400 1.1350 0.5300 1.3750 ;
      RECT 0.4400 1.0450 0.7950 1.1350 ;
      RECT 0.4400 0.8400 0.5300 1.0450 ;
      RECT 0.3000 0.7500 0.5300 0.8400 ;
      RECT 1.2050 1.3100 1.2950 1.8700 ;
      RECT 1.2050 0.4200 1.2950 0.9000 ;
      RECT 0.9150 1.1350 1.0050 1.5250 ;
      RECT 0.9150 1.0450 1.3450 1.1350 ;
      RECT 0.9150 0.7100 1.0050 1.0450 ;
      RECT 1.4650 1.1050 1.8950 1.1950 ;
      RECT 1.4650 1.1950 1.5550 1.5250 ;
      RECT 1.4650 0.7100 1.5550 1.1050 ;
  END
END DLY4_X0P5M_A12TH

MACRO DFFNQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3500 0.3200 0.4500 0.4100 ;
        RECT 0.8700 0.3200 0.9700 0.4200 ;
        RECT 3.9500 0.3200 4.0500 0.5150 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.4650 3.5500 1.6400 ;
        RECT 3.3400 1.2500 3.5500 1.4650 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5200 1.0500 3.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END CKN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9250 0.9500 1.5250 ;
        RECT 0.6100 1.5250 0.9500 1.6250 ;
        RECT 0.5550 0.8250 0.9500 0.9250 ;
        RECT 0.6100 1.6250 0.7100 1.9350 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 2.0950 1.9650 2.1950 2.0800 ;
        RECT 3.9500 1.9500 4.0500 2.0800 ;
        RECT 0.8350 1.8200 1.0050 2.0800 ;
        RECT 0.3400 1.5900 0.4300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.3350 0.6500 1.4250 ;
      RECT 0.5600 1.0400 0.6500 1.3350 ;
      RECT 0.0750 1.4250 0.1700 1.7200 ;
      RECT 0.0750 0.5450 0.1700 1.3350 ;
      RECT 1.4200 1.6750 1.5100 1.7950 ;
      RECT 1.0850 1.5850 1.5100 1.6750 ;
      RECT 1.0850 0.7050 1.1750 1.5850 ;
      RECT 0.2600 0.6150 1.4950 0.7050 ;
      RECT 1.4050 0.4950 1.4950 0.6150 ;
      RECT 0.2600 0.7050 0.3550 1.2150 ;
      RECT 1.7950 1.5950 1.9850 1.6950 ;
      RECT 1.7950 1.4450 1.8850 1.5950 ;
      RECT 1.7950 1.3550 2.4050 1.4450 ;
      RECT 2.3150 1.2350 2.4050 1.3550 ;
      RECT 1.7950 0.7800 1.8850 1.3550 ;
      RECT 1.7950 0.6900 1.9850 0.7800 ;
      RECT 2.5950 1.6050 2.8300 1.6950 ;
      RECT 2.5950 1.1100 2.6850 1.6050 ;
      RECT 2.0100 1.0200 2.6850 1.1100 ;
      RECT 2.0100 1.1100 2.1000 1.2350 ;
      RECT 2.5950 0.7750 2.6850 1.0200 ;
      RECT 2.5950 0.6850 2.8650 0.7750 ;
      RECT 3.1200 1.6000 3.2900 1.6900 ;
      RECT 3.1600 0.6750 3.2500 1.6000 ;
      RECT 2.9550 1.8750 3.7550 1.8900 ;
      RECT 1.6150 1.8000 3.7550 1.8750 ;
      RECT 3.6600 1.7150 3.7550 1.8000 ;
      RECT 3.6600 1.6050 4.1500 1.7150 ;
      RECT 4.0600 0.8950 4.1500 1.6050 ;
      RECT 3.7550 0.8050 4.1500 0.8950 ;
      RECT 1.6150 1.7850 3.0300 1.8000 ;
      RECT 2.9400 1.5150 3.0300 1.7850 ;
      RECT 1.6150 1.4950 1.7050 1.7850 ;
      RECT 2.7750 1.4250 3.0300 1.5150 ;
      RECT 1.2900 1.4050 1.7050 1.4950 ;
      RECT 2.7750 0.8900 2.8650 1.4250 ;
      RECT 1.6150 1.0850 1.7050 1.4050 ;
      RECT 1.5100 0.9950 1.7050 1.0850 ;
      RECT 4.1550 1.8650 4.3450 1.9550 ;
      RECT 4.2550 0.6950 4.3450 1.8650 ;
      RECT 3.3950 0.6050 4.3450 0.6950 ;
      RECT 4.2150 0.4100 4.3450 0.6050 ;
      RECT 3.3950 0.5700 3.4850 0.6050 ;
      RECT 1.6150 0.4800 3.4850 0.5700 ;
      RECT 1.6150 0.5700 1.7050 0.8150 ;
      RECT 2.9550 0.5700 3.0450 1.3150 ;
      RECT 1.2900 0.8150 1.7050 0.9050 ;
      RECT 1.2900 0.9050 1.3950 1.2750 ;
  END
END DFFNQ_X2M_A12TH

MACRO DFFNQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.5600 ;
        RECT 0.8550 0.3200 0.9550 0.4650 ;
        RECT 1.5950 0.3200 1.6850 0.6000 ;
    END
  END VSS

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2600 0.9500 1.4350 ;
        RECT 0.8500 1.0500 1.0600 1.2600 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CKN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1250 1.0100 4.3500 1.2200 ;
        RECT 4.2500 1.2200 4.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0588 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0750 1.4500 0.6950 1.5500 ;
        RECT 0.0750 1.5500 0.1750 1.7200 ;
        RECT 0.5950 1.5500 0.6950 1.8800 ;
        RECT 0.0750 0.7800 0.1700 1.4500 ;
        RECT 0.0750 0.6800 0.6950 0.7800 ;
        RECT 0.0750 0.5400 0.1750 0.6800 ;
        RECT 0.5950 0.4100 0.6950 0.6800 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 2.8050 2.0100 3.0150 2.0800 ;
        RECT 0.3000 1.8950 0.4700 2.0800 ;
        RECT 0.8200 1.8950 0.9900 2.0800 ;
        RECT 1.5350 1.7750 1.7450 2.0800 ;
        RECT 4.3050 1.7400 4.4050 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.3350 0.7200 1.7600 0.8100 ;
      RECT 1.6700 0.8100 1.7600 0.9300 ;
      RECT 0.2900 1.0800 0.7200 1.1700 ;
      RECT 0.6300 0.9600 0.7200 1.0800 ;
      RECT 0.6300 0.8700 1.0200 0.9600 ;
      RECT 0.9300 0.6800 1.0200 0.8700 ;
      RECT 0.9300 0.5900 1.4250 0.6800 ;
      RECT 1.3350 0.6800 1.4250 0.7200 ;
      RECT 1.3350 0.4100 1.4250 0.5900 ;
      RECT 1.3350 0.8100 1.4250 1.4700 ;
      RECT 2.1800 1.4100 2.2700 1.7200 ;
      RECT 1.8500 1.3200 2.2700 1.4100 ;
      RECT 1.8500 1.2450 1.9400 1.3200 ;
      RECT 1.5150 1.1400 1.9400 1.2450 ;
      RECT 1.5150 1.0350 1.6050 1.1400 ;
      RECT 1.8500 0.7700 1.9400 1.1400 ;
      RECT 1.8500 0.6800 2.2550 0.7700 ;
      RECT 2.1650 0.5600 2.2550 0.6800 ;
      RECT 2.5800 1.4150 2.7400 1.6250 ;
      RECT 2.6500 1.0550 2.7400 1.4150 ;
      RECT 2.6500 0.9650 3.1250 1.0550 ;
      RECT 2.6500 0.7600 2.7400 0.9650 ;
      RECT 2.5650 0.6600 2.7400 0.7600 ;
      RECT 3.2150 1.6250 3.6550 1.7150 ;
      RECT 3.2150 1.2850 3.3050 1.6250 ;
      RECT 2.8400 1.1950 3.3050 1.2850 ;
      RECT 3.2150 0.7700 3.3050 1.1950 ;
      RECT 3.2150 0.6800 3.6550 0.7700 ;
      RECT 3.9450 0.6600 4.0350 1.6700 ;
      RECT 4.1250 1.5000 4.5400 1.5900 ;
      RECT 4.4500 0.9700 4.5400 1.5000 ;
      RECT 1.1450 1.5500 1.2400 1.5800 ;
      RECT 1.0400 1.4600 1.2400 1.5500 ;
      RECT 1.1500 0.7900 1.2400 1.4600 ;
      RECT 1.8900 1.8100 2.4700 1.8300 ;
      RECT 3.7650 1.5000 3.8550 1.8300 ;
      RECT 1.8900 1.6700 1.9800 1.8100 ;
      RECT 2.3800 1.2300 2.4700 1.8100 ;
      RECT 3.4350 1.4100 3.8550 1.5000 ;
      RECT 1.1450 1.5800 1.9800 1.6700 ;
      RECT 2.0300 1.1400 2.5600 1.2300 ;
      RECT 3.4350 0.8900 3.5250 1.4100 ;
      RECT 2.0300 1.0600 2.1200 1.1400 ;
      RECT 2.4700 1.0600 2.5600 1.1400 ;
      RECT 1.8900 1.8300 4.2150 1.9200 ;
      RECT 4.1250 1.5900 4.2150 1.8300 ;
      RECT 2.3650 0.4800 4.7200 0.5700 ;
      RECT 4.6300 0.5700 4.7200 1.6700 ;
      RECT 3.6450 1.0950 3.8350 1.1850 ;
      RECT 3.7450 0.5700 3.8350 1.0950 ;
      RECT 2.3650 0.5700 2.4550 0.8600 ;
      RECT 2.1300 0.8600 2.4550 0.9500 ;
  END
END DFFNQ_X3M_A12TH

MACRO DFFNRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.9000 ;
        RECT 2.8350 0.3200 2.9250 0.3950 ;
        RECT 4.4700 0.3200 4.6400 0.3950 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 1.4100 4.0400 1.6500 ;
        RECT 3.9400 0.7050 4.0400 1.4100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9400 1.7500 1.3600 ;
    END
    ANTENNAGATEAREA 0.0669 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 1.1750 2.0250 1.2650 2.0800 ;
        RECT 3.0350 1.9400 3.1250 2.0800 ;
        RECT 0.0800 1.6900 0.1700 2.0800 ;
        RECT 4.5000 1.3500 4.6000 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9800 4.7050 1.1900 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.2850 1.6250 0.4700 1.7150 ;
      RECT 0.2850 0.9400 0.3750 1.6250 ;
      RECT 0.2850 0.8500 0.4300 0.9400 ;
      RECT 0.3400 0.5300 0.4300 0.8500 ;
      RECT 0.5600 1.6150 0.8000 1.7050 ;
      RECT 0.7100 1.1900 0.8000 1.6150 ;
      RECT 0.7100 1.1000 1.3600 1.1900 ;
      RECT 1.2600 0.9700 1.3600 1.1000 ;
      RECT 0.7100 0.6900 0.8000 1.1000 ;
      RECT 0.9500 1.5950 1.9700 1.6850 ;
      RECT 1.8800 0.8500 1.9700 1.5950 ;
      RECT 1.4900 0.7600 1.9700 0.8500 ;
      RECT 0.9500 1.3000 1.0400 1.5950 ;
      RECT 2.0950 1.5950 2.2850 1.6850 ;
      RECT 2.1950 0.8000 2.2850 1.5950 ;
      RECT 2.1950 0.7100 3.2950 0.8000 ;
      RECT 3.0550 0.8000 3.1450 1.1400 ;
      RECT 3.0550 1.1400 3.3650 1.2300 ;
      RECT 2.6600 1.5500 3.5450 1.6400 ;
      RECT 3.4550 1.1900 3.5450 1.5500 ;
      RECT 2.6600 1.0600 2.7500 1.5500 ;
      RECT 3.4550 1.0200 3.8250 1.1900 ;
      RECT 3.4550 0.9000 3.5450 1.0200 ;
      RECT 3.3950 0.7300 3.5450 0.9000 ;
      RECT 0.9250 1.8300 4.2800 1.8400 ;
      RECT 2.4250 1.7500 4.2800 1.8300 ;
      RECT 4.1900 0.6850 4.2800 1.7500 ;
      RECT 0.6450 1.8950 2.5150 1.9200 ;
      RECT 0.9250 1.8400 2.5150 1.8950 ;
      RECT 2.4250 0.9100 2.5150 1.7500 ;
      RECT 0.6450 1.9200 1.0150 1.9850 ;
      RECT 0.5200 0.4850 4.9200 0.5750 ;
      RECT 4.8300 0.5750 4.9200 1.5150 ;
      RECT 0.4750 1.3250 0.6100 1.4950 ;
      RECT 0.5200 0.5750 0.6100 1.3250 ;
  END
END DFFNRPQ_X1M_A12TH

MACRO DFFNRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8450 ;
        RECT 4.8700 0.3200 5.0400 0.3950 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9150 4.3500 1.2900 ;
        RECT 4.1350 1.2900 4.3500 1.3900 ;
        RECT 4.1350 0.8150 4.3500 0.9150 ;
        RECT 4.1350 1.3900 4.2350 1.6600 ;
        RECT 4.1350 0.7050 4.2350 0.8150 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4600 1.0500 1.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 1.2750 2.0250 1.3650 2.0800 ;
        RECT 3.1950 1.9400 3.3650 2.0800 ;
        RECT 0.0800 1.7500 0.1700 2.0800 ;
        RECT 4.9000 1.3800 5.0000 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.9950 5.0750 1.2050 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.2850 1.6400 0.4700 1.7300 ;
      RECT 0.2850 0.9650 0.3750 1.6400 ;
      RECT 0.2850 0.8750 0.4300 0.9650 ;
      RECT 0.3400 0.5350 0.4300 0.8750 ;
      RECT 0.5600 1.6150 0.8150 1.7050 ;
      RECT 0.7250 1.1900 0.8150 1.6150 ;
      RECT 0.7250 1.1000 1.3600 1.1900 ;
      RECT 1.2700 0.9700 1.3600 1.1000 ;
      RECT 0.7250 0.6650 0.8150 1.1000 ;
      RECT 1.0200 1.5950 1.9000 1.6850 ;
      RECT 1.8100 1.4550 1.9000 1.5950 ;
      RECT 1.8100 1.3650 2.0800 1.4550 ;
      RECT 1.9900 1.1000 2.0800 1.3650 ;
      RECT 1.9900 1.0100 2.4850 1.1000 ;
      RECT 2.3950 0.9350 2.4850 1.0100 ;
      RECT 1.9900 0.8500 2.0800 1.0100 ;
      RECT 2.3950 0.8450 2.5650 0.9350 ;
      RECT 1.4900 0.7600 2.0800 0.8500 ;
      RECT 1.0200 1.3000 1.1100 1.5950 ;
      RECT 2.0300 1.5950 2.7850 1.6850 ;
      RECT 2.6950 0.8000 2.7850 1.5950 ;
      RECT 2.6950 0.7550 3.5450 0.8000 ;
      RECT 3.4550 0.8000 3.5450 1.0100 ;
      RECT 2.1800 0.7100 3.5450 0.7550 ;
      RECT 3.4550 1.0100 3.6100 1.1800 ;
      RECT 2.1800 0.7550 2.2700 0.9000 ;
      RECT 2.1800 0.6650 2.8100 0.7100 ;
      RECT 3.6250 1.3600 3.7150 1.6400 ;
      RECT 3.1700 1.2700 3.8150 1.3600 ;
      RECT 3.7250 1.1700 3.8150 1.2700 ;
      RECT 3.1700 0.9150 3.2600 1.2700 ;
      RECT 3.7250 1.0800 3.9550 1.1700 ;
      RECT 3.7250 0.8450 3.8150 1.0800 ;
      RECT 3.6350 0.7550 3.8150 0.8450 ;
      RECT 0.9250 1.8300 4.6800 1.8400 ;
      RECT 2.9250 1.7500 4.6800 1.8300 ;
      RECT 4.5900 0.7250 4.6800 1.7500 ;
      RECT 0.6950 1.8950 3.0150 1.9200 ;
      RECT 0.9250 1.8400 3.0150 1.8950 ;
      RECT 2.9250 0.9300 3.0150 1.7500 ;
      RECT 0.6950 1.9200 1.0150 1.9850 ;
      RECT 0.5200 0.4850 5.3200 0.5750 ;
      RECT 5.2300 0.5750 5.3200 1.5000 ;
      RECT 0.4750 1.3250 0.6100 1.5050 ;
      RECT 0.5200 0.5750 0.6100 1.3250 ;
      RECT 0.7400 0.4700 0.9500 0.4850 ;
  END
END DFFNRPQ_X2M_A12TH

MACRO DFFNRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7500 ;
        RECT 5.1050 0.3200 5.2750 0.3950 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.3900 4.1750 1.6600 ;
        RECT 4.0500 1.2900 4.6900 1.3900 ;
        RECT 4.6000 1.3900 4.6900 1.6600 ;
        RECT 4.5900 0.9150 4.6900 1.2900 ;
        RECT 4.0750 0.8150 4.6900 0.9150 ;
        RECT 4.6000 0.7250 4.6900 0.8150 ;
        RECT 4.0750 0.7050 4.1750 0.8150 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4600 1.0400 1.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 1.2900 2.0100 1.3800 2.0800 ;
        RECT 3.1900 1.9900 3.2900 2.0800 ;
        RECT 3.8150 1.9900 3.9150 2.0800 ;
        RECT 4.3350 1.9900 4.4350 2.0800 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 5.1400 1.4500 5.2400 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1050 1.0100 5.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0396 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.2850 1.6400 0.4700 1.7300 ;
      RECT 0.2850 0.9700 0.3750 1.6400 ;
      RECT 0.2850 0.8800 0.4300 0.9700 ;
      RECT 0.3400 0.5800 0.4300 0.8800 ;
      RECT 0.5600 1.6150 0.8150 1.7050 ;
      RECT 0.7250 1.1450 0.8150 1.6150 ;
      RECT 0.7250 1.0550 1.3600 1.1450 ;
      RECT 1.2700 0.9350 1.3600 1.0550 ;
      RECT 0.7250 0.6900 0.8150 1.0550 ;
      RECT 1.0200 1.5950 1.9200 1.6850 ;
      RECT 1.8300 1.4550 1.9200 1.5950 ;
      RECT 1.8300 1.3650 2.0800 1.4550 ;
      RECT 1.9900 1.1000 2.0800 1.3650 ;
      RECT 1.9900 1.0100 2.4850 1.1000 ;
      RECT 2.3950 0.9350 2.4850 1.0100 ;
      RECT 1.9900 0.8500 2.0800 1.0100 ;
      RECT 2.3950 0.8450 2.5800 0.9350 ;
      RECT 1.4900 0.7600 2.0800 0.8500 ;
      RECT 1.0200 1.2600 1.1100 1.5950 ;
      RECT 2.0300 1.5950 2.7800 1.6850 ;
      RECT 2.6900 0.7550 2.7800 1.5950 ;
      RECT 2.1800 0.6650 3.5050 0.7550 ;
      RECT 2.1800 0.7550 2.2700 0.9000 ;
      RECT 3.4150 0.7550 3.5050 0.9550 ;
      RECT 3.4150 0.9550 3.5700 1.1450 ;
      RECT 3.6850 1.0800 4.3450 1.1700 ;
      RECT 3.5850 1.3600 3.6750 1.6400 ;
      RECT 3.1200 1.2700 3.7750 1.3600 ;
      RECT 3.6850 1.1700 3.7750 1.2700 ;
      RECT 3.1200 0.8950 3.2100 1.2700 ;
      RECT 3.6850 0.8450 3.7750 1.0800 ;
      RECT 3.5950 0.7550 3.7750 0.8450 ;
      RECT 0.9250 1.8300 4.9200 1.8400 ;
      RECT 2.8850 1.7500 4.9200 1.8300 ;
      RECT 4.8300 0.7300 4.9200 1.7500 ;
      RECT 0.6950 1.8950 2.9750 1.9200 ;
      RECT 0.9250 1.8400 2.9750 1.8950 ;
      RECT 2.8850 0.9100 2.9750 1.7500 ;
      RECT 0.6950 1.9200 1.0150 1.9850 ;
      RECT 5.4300 1.3900 5.5200 1.5250 ;
      RECT 5.4300 1.3000 5.5450 1.3900 ;
      RECT 5.4550 0.9000 5.5450 1.3000 ;
      RECT 5.4300 0.8100 5.5450 0.9000 ;
      RECT 5.4300 0.5750 5.5200 0.8100 ;
      RECT 0.5200 0.4850 5.5200 0.5750 ;
      RECT 2.4300 0.4500 2.6400 0.4850 ;
      RECT 0.5200 0.5750 0.6100 1.3250 ;
      RECT 0.7400 0.4600 0.9500 0.4850 ;
      RECT 0.4750 1.3250 0.6100 1.5050 ;
  END
END DFFNRPQ_X3M_A12TH

MACRO DFFNSQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7800 ;
        RECT 1.3500 0.3200 1.4500 0.7500 ;
        RECT 2.9650 0.3200 3.1750 0.5350 ;
        RECT 3.5600 0.3200 3.7700 0.4600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 1.5650 2.0400 1.7750 2.0800 ;
        RECT 0.0750 1.7000 0.1750 2.0800 ;
        RECT 4.4650 1.3850 4.5650 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 1.3850 3.9750 1.6700 ;
        RECT 3.8750 0.7850 3.9750 1.3850 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7950 4.5500 1.1050 ;
        RECT 4.4500 1.1050 4.6500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END CKN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.5150 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.4500 1.8000 1.5500 ;
        RECT 1.7000 1.1750 1.8000 1.4500 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END SN
  OBS
    LAYER M1 ;
      RECT 0.6700 1.8300 4.2350 1.9200 ;
      RECT 4.1450 0.7500 4.2350 1.8300 ;
      RECT 2.0150 1.9200 2.2250 1.9900 ;
      RECT 0.6700 1.9200 0.8800 1.9600 ;
      RECT 2.3650 0.6350 4.8750 0.6600 ;
      RECT 4.7850 0.6600 4.8750 1.5350 ;
      RECT 3.3700 0.5700 4.8750 0.6350 ;
      RECT 4.1400 0.5000 4.3500 0.5700 ;
      RECT 2.3350 1.3650 2.4550 1.5500 ;
      RECT 2.3650 0.7250 2.4550 1.3650 ;
      RECT 2.3650 0.5700 2.4550 0.6350 ;
      RECT 1.6050 0.4800 2.4550 0.5700 ;
      RECT 2.0500 0.4350 2.2600 0.4800 ;
      RECT 2.3650 0.6600 3.4600 0.7250 ;
      RECT 1.1050 0.6050 1.1950 0.8650 ;
      RECT 0.5250 0.5150 1.1950 0.6050 ;
      RECT 0.5250 0.6050 0.6150 1.4800 ;
      RECT 1.6050 0.5700 1.6950 0.8650 ;
      RECT 1.1050 0.8650 1.6950 0.9550 ;
      RECT 0.3400 0.6950 0.4300 1.7700 ;
      RECT 0.7450 1.0800 1.5450 1.1700 ;
      RECT 1.4550 1.1700 1.5450 1.2900 ;
      RECT 0.5400 1.5950 0.8350 1.6850 ;
      RECT 0.7450 1.1700 0.8350 1.5950 ;
      RECT 0.7450 0.7500 0.8350 1.0800 ;
      RECT 1.0050 1.6400 1.9900 1.7400 ;
      RECT 1.8900 0.7000 1.9900 1.6400 ;
      RECT 1.0050 1.2900 1.1050 1.6400 ;
      RECT 2.1300 1.6500 3.1300 1.7400 ;
      RECT 3.0400 1.1700 3.1300 1.6500 ;
      RECT 2.1300 0.9100 2.2200 1.6500 ;
      RECT 3.0400 1.0800 3.4950 1.1700 ;
      RECT 2.1300 0.7000 2.2750 0.9100 ;
      RECT 3.2900 1.3600 3.3800 1.7200 ;
      RECT 3.2900 1.2700 3.7450 1.3600 ;
      RECT 3.6550 0.9350 3.7450 1.2700 ;
      RECT 2.5750 0.8450 3.7450 0.9350 ;
      RECT 2.5750 0.9350 2.6650 1.5350 ;
  END
END DFFNSQ_X1M_A12TH

MACRO DFFNSQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8800 ;
        RECT 1.2650 0.3200 1.4350 0.4500 ;
        RECT 4.5700 0.3200 4.6600 0.7400 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.8700 3.9500 1.2900 ;
        RECT 3.7550 1.2900 3.9500 1.3900 ;
        RECT 3.7550 0.6600 3.9500 0.8700 ;
        RECT 3.7550 1.3900 3.8550 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9600 1.7500 1.5100 ;
    END
    ANTENNAGATEAREA 0.075 ;
  END SN

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6350 1.0300 4.7550 1.4100 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END CKN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 2.6100 2.0100 2.7800 2.0800 ;
        RECT 0.0750 1.7000 0.1750 2.0800 ;
        RECT 4.5200 1.5000 4.6200 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0650 0.1600 1.4500 ;
    END
    ANTENNAGATEAREA 0.0474 ;
  END D
  OBS
    LAYER M1 ;
      RECT 2.0650 1.5800 3.0600 1.6700 ;
      RECT 2.0650 1.5250 2.2500 1.5800 ;
      RECT 2.9700 1.1700 3.0600 1.5800 ;
      RECT 2.0650 0.7200 2.1550 1.5250 ;
      RECT 2.9700 1.0800 3.3750 1.1700 ;
      RECT 3.2000 1.3800 3.2900 1.7200 ;
      RECT 3.2000 1.2900 3.6550 1.3800 ;
      RECT 3.5650 0.8000 3.6550 1.2900 ;
      RECT 2.5350 0.7100 3.6550 0.8000 ;
      RECT 2.5350 0.8000 2.6250 1.4050 ;
      RECT 0.6700 1.8300 4.3000 1.9200 ;
      RECT 4.2100 1.6050 4.3000 1.8300 ;
      RECT 4.2100 1.4350 4.3100 1.6050 ;
      RECT 4.2100 0.6800 4.3000 1.4350 ;
      RECT 2.1600 1.9200 2.3700 1.9900 ;
      RECT 4.8300 1.5900 4.9200 1.7200 ;
      RECT 4.8300 1.5000 4.9550 1.5900 ;
      RECT 4.8650 0.9400 4.9550 1.5000 ;
      RECT 4.3900 0.8500 4.9550 0.9400 ;
      RECT 4.8300 0.6300 4.9200 0.8500 ;
      RECT 4.3900 0.5700 4.4800 0.8500 ;
      RECT 0.5350 0.5400 4.4800 0.5700 ;
      RECT 1.5400 0.4800 4.4800 0.5400 ;
      RECT 4.2150 0.4100 4.4800 0.4800 ;
      RECT 2.3450 0.5700 2.4350 1.2500 ;
      RECT 2.2650 1.2500 2.4350 1.3400 ;
      RECT 1.9350 0.4100 2.1450 0.4800 ;
      RECT 0.8200 0.5250 0.9900 0.5400 ;
      RECT 0.5350 0.6300 0.6250 1.2200 ;
      RECT 0.5200 1.2200 0.6250 1.4300 ;
      RECT 0.5350 0.5700 1.6300 0.6300 ;
      RECT 0.3400 0.5100 0.4300 1.8900 ;
      RECT 0.5400 1.5400 0.8350 1.6300 ;
      RECT 0.7450 0.8450 0.8350 1.5400 ;
      RECT 0.7450 0.7550 1.5300 0.8450 ;
      RECT 1.4400 0.8450 1.5300 1.2500 ;
      RECT 1.3200 1.2500 1.5300 1.3400 ;
      RECT 1.0250 1.6500 1.9450 1.7400 ;
      RECT 1.8550 0.7800 1.9450 1.6500 ;
      RECT 1.7300 0.6900 1.9450 0.7800 ;
      RECT 1.0250 1.1800 1.1150 1.6500 ;
  END
END DFFNSQ_X2M_A12TH

MACRO DFFNSQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.9500 ;
        RECT 1.2650 0.3200 1.4350 0.5150 ;
        RECT 3.4950 0.3200 3.5850 0.3600 ;
        RECT 4.9050 0.3200 4.9950 0.7300 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.7500 4.3650 1.2750 ;
        RECT 3.7550 1.2750 4.3650 1.3750 ;
        RECT 3.7550 0.6600 4.3650 0.7500 ;
        RECT 3.7550 1.3750 3.8550 1.7000 ;
        RECT 4.2750 1.3750 4.3650 1.6900 ;
        RECT 3.7550 0.7500 3.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9600 1.7500 1.5100 ;
    END
    ANTENNAGATEAREA 0.0882 ;
  END SN

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8450 1.0100 4.9550 1.4000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END CKN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 0.0750 1.7950 0.1750 2.0800 ;
        RECT 4.8400 1.5000 4.9400 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0650 0.1600 1.4500 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.5400 1.5400 0.8350 1.6300 ;
      RECT 0.7450 0.9400 0.8350 1.5400 ;
      RECT 0.7450 0.8500 1.4250 0.9400 ;
      RECT 1.3350 0.9400 1.4250 1.2650 ;
      RECT 1.3350 1.2650 1.5500 1.3550 ;
      RECT 1.0250 1.6500 1.9450 1.7400 ;
      RECT 1.8550 0.8300 1.9450 1.6500 ;
      RECT 1.7300 0.7400 1.9450 0.8300 ;
      RECT 1.0250 1.1800 1.1150 1.6500 ;
      RECT 2.0650 1.6300 3.0600 1.7200 ;
      RECT 2.0650 1.5250 2.2500 1.6300 ;
      RECT 2.9700 1.1700 3.0600 1.6300 ;
      RECT 2.0650 0.7600 2.1550 1.5250 ;
      RECT 2.9700 1.0800 3.3750 1.1700 ;
      RECT 3.5650 1.0900 4.0100 1.1800 ;
      RECT 3.2000 1.4150 3.2900 1.7150 ;
      RECT 3.2000 1.3250 3.6550 1.4150 ;
      RECT 3.5650 1.1800 3.6550 1.3250 ;
      RECT 3.5650 0.8000 3.6550 1.0900 ;
      RECT 2.5350 0.7100 3.6550 0.8000 ;
      RECT 2.5350 0.8000 2.6250 1.4200 ;
      RECT 0.6700 1.8300 4.6150 1.9200 ;
      RECT 4.5250 0.6900 4.6150 1.8300 ;
      RECT 2.2250 1.9200 2.4350 1.9900 ;
      RECT 5.1650 1.5900 5.2550 1.7200 ;
      RECT 5.1650 1.5000 5.3500 1.5900 ;
      RECT 5.2600 0.9200 5.3500 1.5000 ;
      RECT 4.7050 0.8300 5.3500 0.9200 ;
      RECT 5.1650 0.6600 5.2550 0.8300 ;
      RECT 0.5200 0.6950 0.6100 1.4300 ;
      RECT 4.7050 0.5700 4.7950 0.8300 ;
      RECT 1.5400 0.4800 4.7950 0.5700 ;
      RECT 4.5400 0.4100 4.7950 0.4800 ;
      RECT 2.3450 0.5700 2.4350 1.2700 ;
      RECT 2.1600 0.4100 2.3700 0.4800 ;
      RECT 2.2650 1.2700 2.4350 1.3600 ;
      RECT 1.5400 0.5700 1.6300 0.6050 ;
      RECT 0.5200 0.6050 1.6300 0.6950 ;
      RECT 0.3400 0.5100 0.4300 1.8900 ;
  END
END DFFNSQ_X3M_A12TH

MACRO DFFNSRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7300 ;
        RECT 2.6050 0.3200 3.0150 0.3700 ;
        RECT 5.5350 0.3200 5.6350 0.6900 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 1.0500 3.1500 1.4750 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1900 4.1500 1.4300 ;
        RECT 3.9050 1.0900 4.1500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0588 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 0.0800 1.7150 0.1700 2.0800 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.8600 4.9500 1.2500 ;
        RECT 4.8500 1.2500 5.0700 1.3500 ;
        RECT 4.8500 0.7600 5.1300 0.8600 ;
        RECT 4.9800 1.3500 5.0700 1.7100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4300 1.0100 5.5500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6400 0.4300 1.7650 ;
      RECT 0.5450 1.5900 0.7900 1.6800 ;
      RECT 0.7000 1.1650 0.7900 1.5900 ;
      RECT 0.7000 1.0750 1.7650 1.1650 ;
      RECT 1.6750 1.1650 1.7650 1.4850 ;
      RECT 0.7000 0.6900 0.7900 1.0750 ;
      RECT 1.5700 0.7600 1.6600 0.9500 ;
      RECT 1.5700 0.6700 2.1800 0.7600 ;
      RECT 2.0900 0.7600 2.1800 0.9400 ;
      RECT 1.0100 1.6200 2.4450 1.7100 ;
      RECT 1.0100 1.2850 1.1000 1.6200 ;
      RECT 2.3400 1.1450 2.4450 1.6200 ;
      RECT 1.8900 1.0550 2.4450 1.1450 ;
      RECT 1.8900 0.9550 1.9800 1.0550 ;
      RECT 2.3550 0.6950 2.4450 1.0550 ;
      RECT 1.7700 0.8650 1.9800 0.9550 ;
      RECT 3.4300 0.6900 4.3850 0.7800 ;
      RECT 4.2950 0.7800 4.3850 1.3250 ;
      RECT 2.6300 1.6450 3.5200 1.7350 ;
      RECT 3.4300 0.7800 3.5200 1.6450 ;
      RECT 2.6300 0.6950 2.7200 1.6450 ;
      RECT 3.8100 1.6400 4.7400 1.7300 ;
      RECT 4.6500 0.7750 4.7400 1.6400 ;
      RECT 4.4750 0.6850 4.7400 0.7750 ;
      RECT 3.8100 1.3300 3.9000 1.6400 ;
      RECT 5.2300 0.8100 5.7550 0.9000 ;
      RECT 5.2300 0.9000 5.3200 1.6750 ;
      RECT 5.2300 0.5700 5.3200 0.8100 ;
      RECT 0.5200 0.4800 5.3200 0.5700 ;
      RECT 3.2400 0.5700 3.3300 1.5350 ;
      RECT 0.5200 0.5700 0.6100 1.4750 ;
      RECT 0.7000 1.8300 5.9350 1.9200 ;
      RECT 5.7950 1.4850 5.9350 1.8300 ;
      RECT 5.8450 0.6700 5.9350 1.4850 ;
      RECT 5.7800 0.4800 5.9350 0.6700 ;
      RECT 3.6300 0.8900 3.7200 1.8300 ;
  END
END DFFNSRPQ_X1M_A12TH

MACRO DFFNSRPQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7600 ;
        RECT 2.7950 0.3200 3.0050 0.3500 ;
        RECT 5.7250 0.3200 5.8150 0.7400 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.2700 2.9500 1.3950 ;
        RECT 2.8500 1.1000 3.1250 1.2700 ;
    END
    ANTENNAGATEAREA 0.0834 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1500 4.1500 1.3900 ;
        RECT 3.8950 1.0500 4.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0714 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.2900 5.0450 1.6600 ;
        RECT 4.8500 0.8600 4.9500 1.2900 ;
        RECT 4.8500 0.7600 5.1050 0.8600 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 1.1700 2.0450 1.3800 2.0800 ;
        RECT 1.9700 2.0450 2.1800 2.0800 ;
        RECT 4.6550 2.0400 4.8250 2.0800 ;
        RECT 4.1900 2.0350 4.3600 2.0800 ;
        RECT 0.0750 1.5500 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9300 0.1600 1.3150 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 1.0400 5.7500 1.4600 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.3400 0.5950 0.4300 1.7200 ;
      RECT 0.5450 1.6900 0.8250 1.7800 ;
      RECT 0.7350 1.1650 0.8250 1.6900 ;
      RECT 0.7350 1.0750 1.7800 1.1650 ;
      RECT 1.6900 1.1650 1.7800 1.2900 ;
      RECT 0.7350 0.6600 0.8250 1.0750 ;
      RECT 1.5700 0.7500 1.6600 0.8700 ;
      RECT 1.5700 0.6600 2.2400 0.7500 ;
      RECT 1.0500 1.5700 1.9750 1.6600 ;
      RECT 1.0500 1.2650 1.1400 1.5700 ;
      RECT 1.8850 0.9300 1.9750 1.5700 ;
      RECT 1.7700 0.8400 2.4600 0.9300 ;
      RECT 2.2750 0.9300 2.3650 1.6350 ;
      RECT 2.3700 0.7200 2.4600 0.8400 ;
      RECT 3.4050 0.6600 4.3850 0.7500 ;
      RECT 4.2950 0.7500 4.3850 1.3450 ;
      RECT 2.5350 1.6450 3.4950 1.7350 ;
      RECT 3.4050 0.7500 3.4950 1.6450 ;
      RECT 2.5350 1.1400 2.6250 1.6450 ;
      RECT 2.5350 1.0500 2.7200 1.1400 ;
      RECT 2.6300 0.7450 2.7200 1.0500 ;
      RECT 3.7950 1.6400 4.6850 1.7300 ;
      RECT 4.5950 0.9250 4.6850 1.6400 ;
      RECT 4.4750 0.7550 4.6850 0.9250 ;
      RECT 3.7950 1.3000 3.8850 1.6400 ;
      RECT 5.4200 0.8300 5.9600 0.9200 ;
      RECT 5.4200 0.9200 5.5100 1.5500 ;
      RECT 5.4200 0.5700 5.5100 0.8300 ;
      RECT 0.5200 0.4800 5.5100 0.5700 ;
      RECT 3.2150 0.5700 3.3050 1.5350 ;
      RECT 0.5200 0.5700 0.6100 1.4700 ;
      RECT 0.7300 1.8950 6.1400 1.9200 ;
      RECT 0.9250 1.8300 6.1400 1.8950 ;
      RECT 6.0500 1.5400 6.1400 1.8300 ;
      RECT 5.9900 1.3300 6.1400 1.5400 ;
      RECT 6.0500 0.7300 6.1400 1.3300 ;
      RECT 6.0000 0.5400 6.1400 0.7300 ;
      RECT 3.6050 0.8650 3.6950 1.8300 ;
      RECT 0.7300 1.9200 1.0150 1.9850 ;
  END
END DFFNSRPQ_X2M_A12TH

MACRO DFFNSRPQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8800 ;
        RECT 2.8400 0.3200 3.0100 0.3800 ;
        RECT 4.6800 0.3200 4.8850 0.3750 ;
        RECT 5.1950 0.3200 5.4050 0.3750 ;
        RECT 6.1150 0.3200 6.2050 0.7300 ;
    END
  END VSS

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.1350 3.1250 1.3050 ;
        RECT 2.8500 1.3050 2.9500 1.4300 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END SN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1500 4.1500 1.3950 ;
        RECT 3.8500 1.0500 4.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9950 1.2500 5.6500 1.3500 ;
        RECT 4.9950 1.3500 5.0950 1.7100 ;
        RECT 5.5200 1.3500 5.6500 1.7100 ;
        RECT 5.4500 0.9500 5.5500 1.2500 ;
        RECT 4.9950 0.8500 5.6700 0.9500 ;
        RECT 4.9950 0.7400 5.0950 0.8500 ;
    END
    ANTENNADIFFAREA 0.595725 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 4.7000 2.0400 4.8700 2.0800 ;
        RECT 1.9500 2.0350 2.1600 2.0800 ;
        RECT 4.1900 2.0350 4.3600 2.0800 ;
        RECT 1.1950 2.0200 1.4050 2.0800 ;
        RECT 0.0800 1.6950 0.1700 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.4650 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END D

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0300 1.0500 6.1500 1.4600 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END CKN
  OBS
    LAYER M1 ;
      RECT 0.3400 0.7600 0.4300 1.9750 ;
      RECT 0.5450 1.5900 0.8250 1.6800 ;
      RECT 0.7350 1.1650 0.8250 1.5900 ;
      RECT 0.7350 1.0750 1.7600 1.1650 ;
      RECT 1.6700 1.1650 1.7600 1.2900 ;
      RECT 0.7350 0.6600 0.8250 1.0750 ;
      RECT 1.5100 0.6600 2.2400 0.7500 ;
      RECT 1.0350 1.5700 1.9750 1.6600 ;
      RECT 1.0350 1.2650 1.1250 1.5700 ;
      RECT 1.8850 0.9300 1.9750 1.5700 ;
      RECT 1.7700 0.8400 2.4600 0.9300 ;
      RECT 2.2750 0.9300 2.3650 1.7250 ;
      RECT 2.3700 0.6650 2.4600 0.8400 ;
      RECT 3.4050 0.6600 4.4000 0.7500 ;
      RECT 4.3100 0.7500 4.4000 1.2300 ;
      RECT 2.5350 1.6450 3.4950 1.7350 ;
      RECT 3.4050 0.7500 3.4950 1.6450 ;
      RECT 2.5350 1.1400 2.6250 1.6450 ;
      RECT 2.5350 1.0500 2.7200 1.1400 ;
      RECT 2.6300 0.6650 2.7200 1.0500 ;
      RECT 4.4900 1.0600 5.3350 1.1500 ;
      RECT 3.7950 1.6400 4.5800 1.7300 ;
      RECT 4.4900 1.1500 4.5800 1.6400 ;
      RECT 4.4900 0.7500 4.5800 1.0600 ;
      RECT 3.7950 1.3000 3.8850 1.6400 ;
      RECT 5.8000 0.8300 6.3350 0.9200 ;
      RECT 0.5200 0.4800 5.8900 0.5700 ;
      RECT 5.8000 0.5700 5.8900 0.8300 ;
      RECT 5.8000 0.9200 5.8900 1.6300 ;
      RECT 3.2150 1.0250 3.3050 1.5350 ;
      RECT 2.8100 0.9350 3.3050 1.0250 ;
      RECT 3.2150 0.5700 3.3050 0.9350 ;
      RECT 0.5200 0.5700 0.6100 1.4750 ;
      RECT 0.7300 1.8300 6.5500 1.9200 ;
      RECT 6.4100 1.4800 6.5500 1.8300 ;
      RECT 6.4600 0.7300 6.5500 1.4800 ;
      RECT 6.4150 0.5200 6.5500 0.7300 ;
      RECT 3.6050 0.8650 3.6950 1.8300 ;
  END
END DFFNSRPQ_X3M_A12TH

MACRO DFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.8500 ;
        RECT 3.6950 0.3200 3.8650 0.7300 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.7750 3.1500 1.6150 ;
        RECT 3.0500 1.6150 3.3250 1.7150 ;
        RECT 3.0500 0.6750 3.3250 0.7750 ;
    END
    ANTENNADIFFAREA 0.14175 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.0550 1.5850 0.2250 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.2400 1.2250 ;
    END
    ANTENNAGATEAREA 0.0192 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8450 1.0550 3.9500 1.4750 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3300 1.5500 0.4450 1.7400 ;
      RECT 0.3300 0.8500 0.4200 1.5500 ;
      RECT 0.3300 0.6400 0.4450 0.8500 ;
      RECT 0.5550 1.5900 0.8400 1.6800 ;
      RECT 0.7500 1.0550 0.8400 1.5900 ;
      RECT 0.7500 0.9650 1.4300 1.0550 ;
      RECT 1.3400 1.0550 1.4300 1.2900 ;
      RECT 0.7500 0.6600 0.8400 0.9650 ;
      RECT 1.0150 1.5800 1.6400 1.6700 ;
      RECT 1.0150 1.1550 1.1050 1.5800 ;
      RECT 1.5500 0.6600 1.6400 1.5800 ;
      RECT 2.4250 1.0850 2.6850 1.1750 ;
      RECT 2.4250 0.8050 2.5150 1.0850 ;
      RECT 1.7500 0.7150 2.5150 0.8050 ;
      RECT 1.7500 0.8050 1.8400 1.7300 ;
      RECT 2.1450 1.5750 2.9200 1.6650 ;
      RECT 2.1450 1.2000 2.2350 1.5750 ;
      RECT 2.8200 0.8050 2.9200 1.5750 ;
      RECT 2.6400 0.7150 2.9200 0.8050 ;
      RECT 0.5500 0.4800 3.5300 0.5700 ;
      RECT 3.4400 0.5700 3.5300 1.7300 ;
      RECT 0.5100 1.3150 0.6400 1.4850 ;
      RECT 0.5500 0.5700 0.6400 1.3150 ;
      RECT 0.7200 1.8200 3.9850 1.9100 ;
      RECT 3.8950 1.6750 3.9850 1.8200 ;
      RECT 3.8950 1.5750 4.1550 1.6750 ;
      RECT 4.0650 0.9550 4.1550 1.5750 ;
      RECT 3.6200 0.8650 4.1550 0.9550 ;
      RECT 4.0650 0.7300 4.1550 0.8650 ;
      RECT 3.9550 0.6400 4.1550 0.7300 ;
      RECT 1.9550 0.9150 2.0450 1.8200 ;
  END
END DFFQN_X0P5M_A12TH

MACRO DFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.8000 ;
        RECT 2.8750 0.3200 3.0550 0.3750 ;
        RECT 3.6950 0.3200 3.8650 0.7300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.0950 1.5250 0.1850 2.0800 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9450 3.1500 1.3800 ;
        RECT 3.0500 1.3800 3.3250 1.4800 ;
        RECT 3.0500 0.8450 3.3250 0.9450 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.2400 1.2250 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8450 1.0550 3.9500 1.4750 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3300 1.5650 0.4450 1.7750 ;
      RECT 0.3300 0.8400 0.4200 1.5650 ;
      RECT 0.3300 0.6100 0.4450 0.8400 ;
      RECT 0.5550 1.5900 0.8400 1.6800 ;
      RECT 0.7500 1.0550 0.8400 1.5900 ;
      RECT 0.7500 0.9650 1.4300 1.0550 ;
      RECT 1.3400 1.0550 1.4300 1.3750 ;
      RECT 0.7500 0.6850 0.8400 0.9650 ;
      RECT 1.0150 1.5800 1.6500 1.6700 ;
      RECT 1.0150 1.1550 1.1050 1.5800 ;
      RECT 1.5600 0.6700 1.6500 1.5800 ;
      RECT 2.3750 1.0850 2.7550 1.1750 ;
      RECT 2.3750 0.8500 2.4650 1.0850 ;
      RECT 1.7700 0.7600 2.4650 0.8500 ;
      RECT 1.7700 0.8500 1.8600 1.7400 ;
      RECT 2.1750 1.5750 2.9450 1.6650 ;
      RECT 2.1750 1.2000 2.2650 1.5750 ;
      RECT 2.8450 0.8500 2.9450 1.5750 ;
      RECT 2.6600 0.7600 2.9450 0.8500 ;
      RECT 0.5500 0.4800 3.5300 0.5700 ;
      RECT 3.4400 0.5700 3.5300 1.7300 ;
      RECT 0.5100 1.3300 0.6400 1.5000 ;
      RECT 0.5500 0.5700 0.6400 1.3300 ;
      RECT 1.6900 0.4200 1.9050 0.4800 ;
      RECT 0.7200 1.8300 3.9850 1.9200 ;
      RECT 3.8950 1.6750 3.9850 1.8300 ;
      RECT 3.8950 1.5850 4.1550 1.6750 ;
      RECT 4.0650 0.9550 4.1550 1.5850 ;
      RECT 3.6200 0.8650 4.1550 0.9550 ;
      RECT 4.0650 0.7300 4.1550 0.8650 ;
      RECT 3.9550 0.6400 4.1550 0.7300 ;
      RECT 1.5900 1.9200 1.7600 1.9900 ;
      RECT 1.9850 0.9400 2.0750 1.8300 ;
  END
END DFFQN_X1M_A12TH

MACRO DFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.5200 ;
        RECT 0.8750 0.3200 1.0450 0.5200 ;
        RECT 2.1550 0.3200 2.5250 0.3800 ;
        RECT 3.9200 0.3200 4.0900 0.5050 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.8550 3.5500 1.2850 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7450 1.6500 4.1650 1.7500 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9300 0.7850 1.3050 ;
        RECT 0.5850 1.3050 0.7850 1.3950 ;
        RECT 0.5950 0.8200 0.7850 0.9300 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 3.5450 2.0000 3.6650 2.0800 ;
        RECT 3.9550 1.8800 4.0550 2.0800 ;
        RECT 0.3900 1.7950 0.4900 2.0800 ;
        RECT 0.9050 1.7950 1.0200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0900 1.4900 1.0800 1.5800 ;
      RECT 0.9900 1.0150 1.0800 1.4900 ;
      RECT 0.0900 0.7500 0.1850 1.4900 ;
      RECT 1.5000 1.6750 1.5950 1.7800 ;
      RECT 1.1700 1.5850 1.5950 1.6750 ;
      RECT 1.1700 0.7000 1.2600 1.5850 ;
      RECT 0.3900 0.6100 1.6250 0.7000 ;
      RECT 1.5300 0.4950 1.6250 0.6100 ;
      RECT 0.3900 0.7000 0.4850 1.2350 ;
      RECT 1.8950 1.5900 2.5150 1.6900 ;
      RECT 2.4100 1.1100 2.5150 1.5900 ;
      RECT 1.8950 0.8100 1.9850 1.5900 ;
      RECT 1.8950 0.7150 2.0850 0.8100 ;
      RECT 2.6700 1.6050 2.9100 1.6950 ;
      RECT 2.6700 0.9900 2.7600 1.6050 ;
      RECT 2.0950 0.9000 2.7600 0.9900 ;
      RECT 2.0950 0.9900 2.1850 1.3450 ;
      RECT 2.6700 0.7750 2.7600 0.9000 ;
      RECT 2.6700 0.6850 2.9400 0.7750 ;
      RECT 3.2300 0.6600 3.3200 1.7200 ;
      RECT 3.4100 1.4550 4.0050 1.5450 ;
      RECT 3.9000 0.7950 4.0050 1.4550 ;
      RECT 1.6850 1.8300 3.5000 1.9200 ;
      RECT 3.4100 1.5450 3.5000 1.8300 ;
      RECT 3.0200 1.5150 3.1100 1.8300 ;
      RECT 1.6850 1.4950 1.7750 1.8300 ;
      RECT 2.8500 1.4250 3.1100 1.5150 ;
      RECT 1.3750 1.4050 1.7750 1.4950 ;
      RECT 2.8500 0.8850 2.9400 1.4250 ;
      RECT 1.6850 1.0900 1.7750 1.4050 ;
      RECT 1.5650 0.9950 1.7750 1.0900 ;
      RECT 4.1650 1.8650 4.3500 1.9550 ;
      RECT 4.2550 0.6850 4.3500 1.8650 ;
      RECT 3.7050 0.5950 4.3500 0.6850 ;
      RECT 4.2200 0.4100 4.3500 0.5950 ;
      RECT 3.7050 0.6850 3.7950 1.2950 ;
      RECT 3.7050 0.5700 3.7950 0.5950 ;
      RECT 1.7150 0.4800 3.7950 0.5700 ;
      RECT 1.7150 0.5700 1.8050 0.8150 ;
      RECT 3.0300 0.5700 3.1200 1.3150 ;
      RECT 1.3550 0.8150 1.8050 0.9050 ;
      RECT 1.3550 0.9050 1.4550 1.2850 ;
  END
END DFFQN_X2M_A12TH

MACRO DFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.3500 0.3200 0.5200 0.5200 ;
        RECT 0.8700 0.3200 1.0400 0.5200 ;
        RECT 1.3650 0.3200 1.4650 0.5200 ;
        RECT 3.8850 0.3200 4.0900 0.3900 ;
        RECT 4.3200 0.3200 4.4900 0.5050 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.8550 3.9500 1.2850 ;
    END
    ANTENNAGATEAREA 0.0642 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1450 1.6500 4.5650 1.7500 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9300 1.1500 1.3050 ;
        RECT 0.5900 1.3050 1.3050 1.3950 ;
        RECT 0.5950 0.9150 1.1500 0.9300 ;
        RECT 0.5950 0.8250 1.3150 0.9150 ;
    END
    ANTENNADIFFAREA 0.5415 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 3.9100 1.9800 4.1000 2.0800 ;
        RECT 4.3550 1.8800 4.4550 2.0800 ;
        RECT 0.3850 1.7950 0.4850 2.0800 ;
        RECT 0.8950 1.7950 1.0100 2.0800 ;
        RECT 1.3700 1.7100 1.4700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0900 1.5050 1.4850 1.5950 ;
      RECT 1.3950 1.0150 1.4850 1.5050 ;
      RECT 0.0900 0.7500 0.1850 1.5050 ;
      RECT 1.9100 1.6750 2.0050 1.7800 ;
      RECT 1.5750 1.5850 2.0050 1.6750 ;
      RECT 1.5750 0.7000 1.6650 1.5850 ;
      RECT 0.3000 0.6100 2.0250 0.7000 ;
      RECT 1.9300 0.4950 2.0250 0.6100 ;
      RECT 0.3000 0.7000 0.3950 1.0550 ;
      RECT 0.3000 1.0550 0.9500 1.1550 ;
      RECT 2.2950 1.5900 2.9150 1.6900 ;
      RECT 2.8100 1.1100 2.9150 1.5900 ;
      RECT 2.2950 0.8100 2.3850 1.5900 ;
      RECT 2.2950 0.7150 2.4850 0.8100 ;
      RECT 3.0700 1.6050 3.3100 1.6950 ;
      RECT 3.0700 0.9900 3.1600 1.6050 ;
      RECT 2.4950 0.9000 3.1600 0.9900 ;
      RECT 2.4950 0.9900 2.5850 1.2050 ;
      RECT 3.0700 0.7700 3.1600 0.9000 ;
      RECT 3.0700 0.6800 3.3400 0.7700 ;
      RECT 3.6300 0.6600 3.7200 1.7100 ;
      RECT 3.8300 1.4500 4.4050 1.5400 ;
      RECT 4.3000 0.7950 4.4050 1.4500 ;
      RECT 2.0950 1.8000 3.9200 1.8900 ;
      RECT 3.8300 1.5400 3.9200 1.8000 ;
      RECT 3.4200 1.5100 3.5100 1.8000 ;
      RECT 2.0950 1.4950 2.1850 1.8000 ;
      RECT 3.2500 1.4200 3.5100 1.5100 ;
      RECT 1.7750 1.4050 2.1850 1.4950 ;
      RECT 3.2500 0.8800 3.3400 1.4200 ;
      RECT 2.0950 1.0900 2.1850 1.4050 ;
      RECT 1.9950 0.9950 2.1850 1.0900 ;
      RECT 4.5650 1.8650 4.7500 1.9550 ;
      RECT 4.6550 0.6850 4.7500 1.8650 ;
      RECT 4.1050 0.5950 4.7500 0.6850 ;
      RECT 4.6200 0.4100 4.7500 0.5950 ;
      RECT 4.1050 0.6850 4.1950 1.2950 ;
      RECT 4.1050 0.5700 4.1950 0.5950 ;
      RECT 2.1150 0.4800 4.1950 0.5700 ;
      RECT 2.1150 0.5700 2.2050 0.8150 ;
      RECT 3.4300 0.5700 3.5200 1.3100 ;
      RECT 1.7850 0.8150 2.2050 0.9050 ;
      RECT 1.7850 0.9050 1.8850 1.2850 ;
  END
END DFFQN_X3M_A12TH

MACRO DFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3250 0.3200 0.4950 0.5250 ;
        RECT 0.8100 0.3200 0.9800 0.4650 ;
        RECT 2.1200 0.3200 2.4900 0.3800 ;
        RECT 3.4250 0.3200 3.7950 0.3700 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.9600 3.3500 1.1300 ;
        RECT 3.2500 1.1300 3.4000 1.3000 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5500 1.6500 3.9750 1.7500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9150 0.9500 1.5400 ;
        RECT 0.6500 1.5400 0.9500 1.6300 ;
        RECT 0.5950 0.8150 0.9500 0.9150 ;
        RECT 0.6500 1.6300 0.7500 1.7300 ;
    END
    ANTENNADIFFAREA 0.1304 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 3.1800 2.0150 3.5500 2.0800 ;
        RECT 2.0850 1.9750 2.4550 2.0800 ;
        RECT 3.7500 1.8800 3.8500 2.0800 ;
        RECT 0.8800 1.7500 0.9800 2.0800 ;
        RECT 0.3800 1.5600 0.4800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.3600 0.7050 1.4500 ;
      RECT 0.6150 1.0450 0.7050 1.3600 ;
      RECT 0.0750 0.7350 0.1700 1.3600 ;
      RECT 1.4100 1.6750 1.5050 1.7750 ;
      RECT 1.0650 1.5850 1.5050 1.6750 ;
      RECT 1.0650 0.7050 1.1550 1.5850 ;
      RECT 0.2600 0.6150 1.5050 0.7050 ;
      RECT 1.4100 0.4950 1.5050 0.6150 ;
      RECT 0.2600 0.7050 0.3550 1.2350 ;
      RECT 1.7750 1.5950 2.3900 1.6900 ;
      RECT 2.2950 1.1100 2.3900 1.5950 ;
      RECT 1.7750 0.7750 1.8650 1.5950 ;
      RECT 1.7750 0.6800 1.9650 0.7750 ;
      RECT 2.4950 1.6050 2.7650 1.6950 ;
      RECT 2.4950 0.9900 2.5850 1.6050 ;
      RECT 1.9700 0.9000 2.5850 0.9900 ;
      RECT 1.9700 0.9900 2.0600 1.4150 ;
      RECT 2.4950 0.7700 2.5850 0.9000 ;
      RECT 2.4950 0.6800 2.7950 0.7700 ;
      RECT 3.0700 1.4750 3.1800 1.6450 ;
      RECT 3.0700 0.6800 3.1600 1.4750 ;
      RECT 3.2700 1.4050 3.8550 1.4950 ;
      RECT 3.7450 0.7250 3.8550 1.4050 ;
      RECT 1.5950 1.7850 3.3600 1.8750 ;
      RECT 3.2700 1.4950 3.3600 1.7850 ;
      RECT 2.8800 1.5150 2.9700 1.7850 ;
      RECT 1.5950 1.4950 1.6850 1.7850 ;
      RECT 2.6750 1.4250 2.9700 1.5150 ;
      RECT 1.2650 1.4050 1.6850 1.4950 ;
      RECT 2.6750 0.8850 2.7650 1.4250 ;
      RECT 1.5950 1.0850 1.6850 1.4050 ;
      RECT 1.4900 0.9950 1.6850 1.0850 ;
      RECT 3.9650 1.8800 4.1550 1.9700 ;
      RECT 4.0650 0.6600 4.1550 1.8800 ;
      RECT 4.0200 0.5700 4.1550 0.6600 ;
      RECT 1.5950 0.4800 4.1200 0.5700 ;
      RECT 4.0200 0.4100 4.1200 0.4800 ;
      RECT 3.5600 0.5700 3.6500 1.2950 ;
      RECT 1.5950 0.5700 1.6850 0.8150 ;
      RECT 2.8850 0.5700 2.9750 1.3150 ;
      RECT 1.2800 0.8150 1.6850 0.9050 ;
      RECT 1.2800 0.9050 1.3800 1.2850 ;
  END
END DFFQ_X0P5M_A12TH

MACRO DFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.5200 ;
        RECT 0.8100 0.3200 0.9800 0.4650 ;
        RECT 2.1200 0.3200 2.4900 0.3800 ;
        RECT 3.4250 0.3200 3.7950 0.3700 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.9600 3.3500 1.1300 ;
        RECT 3.2500 1.1300 3.4000 1.3000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5550 1.6500 3.9750 1.7500 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9100 0.9500 1.5400 ;
        RECT 0.6400 1.5400 0.9500 1.6300 ;
        RECT 0.5950 0.8100 0.9500 0.9100 ;
        RECT 0.6400 1.6300 0.7400 1.9400 ;
    END
    ANTENNADIFFAREA 0.238675 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 2.0850 1.9750 2.4550 2.0800 ;
        RECT 3.7500 1.8800 3.8500 2.0800 ;
        RECT 0.3800 1.7700 0.4800 2.0800 ;
        RECT 0.8900 1.7500 0.9900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.3600 0.7050 1.4500 ;
      RECT 0.6150 1.0450 0.7050 1.3600 ;
      RECT 0.0800 1.4500 0.1700 1.7200 ;
      RECT 0.0800 0.7200 0.1700 1.3600 ;
      RECT 1.4100 1.6750 1.5050 1.7750 ;
      RECT 1.0650 1.5850 1.5050 1.6750 ;
      RECT 1.0650 0.7000 1.1550 1.5850 ;
      RECT 0.2600 0.6100 1.5050 0.7000 ;
      RECT 1.4100 0.5100 1.5050 0.6100 ;
      RECT 0.2600 0.7000 0.3550 1.2350 ;
      RECT 1.7750 1.5950 2.3900 1.6900 ;
      RECT 2.2950 1.1100 2.3900 1.5950 ;
      RECT 1.7750 0.7750 1.8650 1.5950 ;
      RECT 1.7750 0.6800 1.9650 0.7750 ;
      RECT 2.4950 1.6050 2.7650 1.6950 ;
      RECT 2.4950 0.9900 2.5850 1.6050 ;
      RECT 1.9700 0.9000 2.5850 0.9900 ;
      RECT 1.9700 0.9900 2.0600 1.4150 ;
      RECT 2.4950 0.7700 2.5850 0.9000 ;
      RECT 2.4950 0.6800 2.7950 0.7700 ;
      RECT 3.0700 0.6800 3.1600 1.6650 ;
      RECT 3.2700 1.4050 3.8550 1.4950 ;
      RECT 3.7450 0.7250 3.8550 1.4050 ;
      RECT 1.5950 1.7850 3.3600 1.8750 ;
      RECT 3.2700 1.4950 3.3600 1.7850 ;
      RECT 2.8800 1.5150 2.9700 1.7850 ;
      RECT 1.5950 1.4950 1.6850 1.7850 ;
      RECT 2.6750 1.4250 2.9700 1.5150 ;
      RECT 1.2650 1.4050 1.6850 1.4950 ;
      RECT 2.6750 0.8850 2.7650 1.4250 ;
      RECT 1.5950 1.0850 1.6850 1.4050 ;
      RECT 1.4900 0.9950 1.6850 1.0850 ;
      RECT 3.9650 1.8800 4.1550 1.9700 ;
      RECT 4.0650 0.6600 4.1550 1.8800 ;
      RECT 4.0200 0.5700 4.1550 0.6600 ;
      RECT 1.5950 0.4800 4.1200 0.5700 ;
      RECT 4.0200 0.4100 4.1200 0.4800 ;
      RECT 3.5600 0.5700 3.6500 1.2950 ;
      RECT 1.5950 0.5700 1.6850 0.8150 ;
      RECT 2.8850 0.5700 2.9750 1.3150 ;
      RECT 1.2800 0.8150 1.6850 0.9050 ;
      RECT 1.2800 0.9050 1.3800 1.2850 ;
  END
END DFFQ_X1M_A12TH

MACRO DFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.3800 0.3200 0.4800 0.4500 ;
        RECT 0.8750 0.3200 1.0450 0.5250 ;
        RECT 3.9200 0.3200 4.0900 0.4800 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.8550 3.5500 1.2850 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7450 1.6500 4.1650 1.7550 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.9300 0.9500 1.5250 ;
        RECT 0.6400 1.5250 0.9500 1.6150 ;
        RECT 0.5850 0.8300 0.9500 0.9300 ;
        RECT 0.6400 1.6150 0.7400 1.9200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 2.1650 1.9650 2.2700 2.0800 ;
        RECT 3.9500 1.9250 4.0500 2.0800 ;
        RECT 0.9250 1.7700 1.0400 2.0800 ;
        RECT 0.3450 1.6200 0.4450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.3450 0.7050 1.4350 ;
      RECT 0.6150 1.0450 0.7050 1.3450 ;
      RECT 0.0750 1.4350 0.1700 1.7350 ;
      RECT 0.0750 0.5650 0.1700 1.3450 ;
      RECT 1.4850 1.6750 1.5800 1.7750 ;
      RECT 1.1100 1.5850 1.5800 1.6750 ;
      RECT 1.1100 0.7050 1.2000 1.5850 ;
      RECT 0.2600 0.6150 1.5800 0.7050 ;
      RECT 1.4850 0.4950 1.5800 0.6150 ;
      RECT 0.2600 0.7050 0.3550 1.2350 ;
      RECT 1.8500 1.5950 2.5150 1.6900 ;
      RECT 2.4150 1.1100 2.5150 1.5950 ;
      RECT 1.8500 0.8100 1.9400 1.5950 ;
      RECT 1.8500 0.7150 2.0350 0.8100 ;
      RECT 2.6700 1.6050 2.9100 1.6950 ;
      RECT 2.6700 0.9900 2.7600 1.6050 ;
      RECT 2.0650 0.9000 2.7600 0.9900 ;
      RECT 2.0650 0.9900 2.1550 1.4150 ;
      RECT 2.6700 0.7750 2.7600 0.9000 ;
      RECT 2.6700 0.6850 2.9400 0.7750 ;
      RECT 3.2300 0.6600 3.3200 1.6400 ;
      RECT 3.4100 1.4700 3.9950 1.5600 ;
      RECT 3.8850 0.7850 3.9950 1.4700 ;
      RECT 1.6700 1.7850 3.5000 1.8750 ;
      RECT 3.4100 1.5600 3.5000 1.7850 ;
      RECT 3.0200 1.5150 3.1100 1.7850 ;
      RECT 1.6700 1.4950 1.7600 1.7850 ;
      RECT 2.8500 1.4250 3.1100 1.5150 ;
      RECT 1.3250 1.4050 1.7600 1.4950 ;
      RECT 2.8500 0.8850 2.9400 1.4250 ;
      RECT 1.6700 1.0850 1.7600 1.4050 ;
      RECT 1.5650 0.9950 1.7600 1.0850 ;
      RECT 4.1600 1.8650 4.3500 1.9550 ;
      RECT 4.2550 0.6600 4.3500 1.8650 ;
      RECT 3.7050 0.5700 4.3500 0.6600 ;
      RECT 4.2300 0.4100 4.3500 0.5700 ;
      RECT 3.7050 0.6600 3.7950 1.2300 ;
      RECT 1.6700 0.4800 3.7950 0.5700 ;
      RECT 1.6700 0.5700 1.7600 0.8150 ;
      RECT 3.0300 0.5700 3.1200 1.3150 ;
      RECT 1.3550 0.8150 1.7600 0.9050 ;
      RECT 1.3550 0.9050 1.4550 1.2850 ;
  END
END DFFQ_X2M_A12TH

MACRO DFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.3800 0.3200 0.4800 0.4500 ;
        RECT 0.8650 0.3200 1.0350 0.5250 ;
        RECT 4.3150 0.3200 4.4850 0.4650 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.8550 3.9500 1.2850 ;
    END
    ANTENNAGATEAREA 0.0588 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1450 1.6500 4.5650 1.7550 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5850 0.8300 1.3300 0.9300 ;
        RECT 0.5850 0.9300 1.2550 0.9500 ;
        RECT 1.1550 0.9500 1.2550 1.5250 ;
        RECT 0.6400 1.5250 1.2550 1.6150 ;
        RECT 0.6400 1.6150 0.7400 1.9500 ;
        RECT 1.1650 1.6150 1.2550 1.9500 ;
    END
    ANTENNADIFFAREA 0.560025 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 4.3500 1.9900 4.4500 2.0800 ;
        RECT 2.5650 1.9650 2.6700 2.0800 ;
        RECT 0.9000 1.7900 1.0000 2.0800 ;
        RECT 0.3450 1.7700 0.4450 2.0800 ;
        RECT 1.3950 1.5750 1.4850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.3450 0.6600 1.4350 ;
      RECT 0.5700 1.1800 0.6600 1.3450 ;
      RECT 0.5700 1.0900 0.9400 1.1800 ;
      RECT 0.0750 1.4350 0.1700 1.7350 ;
      RECT 0.0750 0.5650 0.1700 1.3450 ;
      RECT 1.9050 1.6750 2.0000 1.8800 ;
      RECT 1.5750 1.5850 2.0000 1.6750 ;
      RECT 1.5750 0.7050 1.6650 1.5850 ;
      RECT 0.2600 0.6150 2.0000 0.7050 ;
      RECT 1.9050 0.4350 2.0000 0.6150 ;
      RECT 0.2600 0.7050 0.3550 1.2350 ;
      RECT 2.2700 1.5950 2.9150 1.6900 ;
      RECT 2.8150 1.1100 2.9150 1.5950 ;
      RECT 2.2700 0.7750 2.3600 1.5950 ;
      RECT 2.2700 0.6800 2.4550 0.7750 ;
      RECT 3.0700 1.6050 3.3100 1.6950 ;
      RECT 3.0700 0.9900 3.1600 1.6050 ;
      RECT 2.4650 0.9000 3.1600 0.9900 ;
      RECT 2.4650 0.9900 2.5550 1.3700 ;
      RECT 3.0700 0.7750 3.1600 0.9000 ;
      RECT 3.0700 0.6850 3.3400 0.7750 ;
      RECT 3.6300 0.6600 3.7200 1.6150 ;
      RECT 3.8100 1.4700 4.3950 1.5600 ;
      RECT 4.2850 0.7900 4.3950 1.4700 ;
      RECT 2.0900 1.7850 3.9000 1.8750 ;
      RECT 3.8100 1.5600 3.9000 1.7850 ;
      RECT 3.4200 1.5150 3.5100 1.7850 ;
      RECT 2.0900 1.4950 2.1800 1.7850 ;
      RECT 3.2500 1.4250 3.5100 1.5150 ;
      RECT 1.7750 1.4050 2.1800 1.4950 ;
      RECT 3.2500 0.8850 3.3400 1.4250 ;
      RECT 2.0900 1.0850 2.1800 1.4050 ;
      RECT 1.9850 0.9950 2.1800 1.0850 ;
      RECT 4.5600 1.9000 4.7500 1.9900 ;
      RECT 4.6550 0.6600 4.7500 1.9000 ;
      RECT 4.1050 0.5700 4.7500 0.6600 ;
      RECT 4.6300 0.4100 4.7500 0.5700 ;
      RECT 4.1050 0.6600 4.1950 1.2700 ;
      RECT 2.0900 0.4800 4.1950 0.5700 ;
      RECT 3.4300 0.5700 3.5200 1.3150 ;
      RECT 2.0900 0.5700 2.1800 0.8150 ;
      RECT 1.7800 0.8150 2.1800 0.9050 ;
      RECT 1.7800 0.9050 1.8700 1.2850 ;
  END
END DFFQ_X3M_A12TH

MACRO DFFQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.5900 0.3200 0.7000 0.4500 ;
        RECT 1.1100 0.3200 1.2150 0.4500 ;
        RECT 1.6000 0.3200 1.7700 0.5250 ;
        RECT 4.7150 0.3200 4.8900 0.4200 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.8550 4.3500 1.2850 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5450 1.6500 4.9650 1.7500 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8000 0.8300 1.7500 0.9500 ;
        RECT 1.6500 0.9500 1.7500 1.5250 ;
        RECT 0.8550 1.5250 1.7500 1.6150 ;
        RECT 0.8550 1.6150 0.9550 1.9450 ;
        RECT 1.3750 1.6150 1.4750 1.9450 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 2.9650 1.9900 3.0700 2.0800 ;
        RECT 4.7500 1.8400 4.8500 2.0800 ;
        RECT 1.1150 1.7900 1.2150 2.0800 ;
        RECT 1.6350 1.7900 1.7350 2.0800 ;
        RECT 0.5950 1.5400 0.6950 2.0800 ;
        RECT 0.0750 1.5350 0.1750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7450 1.0900 1.5150 1.1800 ;
      RECT 0.1900 1.3450 0.8350 1.4350 ;
      RECT 0.7450 1.1800 0.8350 1.3450 ;
      RECT 0.3350 1.4350 0.4350 1.7650 ;
      RECT 0.1900 0.8650 0.2850 1.3450 ;
      RECT 0.1900 0.7750 0.4350 0.8650 ;
      RECT 0.3350 0.4700 0.4350 0.7750 ;
      RECT 2.3050 1.6950 2.4000 1.9900 ;
      RECT 1.9500 1.6050 2.4000 1.6950 ;
      RECT 1.9500 0.7050 2.0400 1.6050 ;
      RECT 0.5400 0.6150 2.4000 0.7050 ;
      RECT 2.3050 0.4350 2.4000 0.6150 ;
      RECT 0.5400 0.7050 0.6350 1.0950 ;
      RECT 0.3750 1.0950 0.6350 1.1850 ;
      RECT 2.6700 1.5950 3.3150 1.6900 ;
      RECT 3.2150 1.1100 3.3150 1.5950 ;
      RECT 2.6700 0.8100 2.7600 1.5950 ;
      RECT 2.6700 0.7150 2.8550 0.8100 ;
      RECT 3.4700 1.6050 3.7100 1.6950 ;
      RECT 3.4700 0.9900 3.5600 1.6050 ;
      RECT 2.8650 0.9000 3.5600 0.9900 ;
      RECT 2.8650 0.9900 2.9550 1.3000 ;
      RECT 3.4700 0.7750 3.5600 0.9000 ;
      RECT 3.4700 0.6850 3.7400 0.7750 ;
      RECT 4.0300 0.6600 4.1200 1.6250 ;
      RECT 4.2100 1.4150 4.7950 1.5050 ;
      RECT 4.6850 0.7900 4.7950 1.4150 ;
      RECT 2.4900 1.7850 4.3000 1.8750 ;
      RECT 4.2100 1.5050 4.3000 1.7850 ;
      RECT 3.8200 1.5150 3.9100 1.7850 ;
      RECT 2.4900 1.4950 2.5800 1.7850 ;
      RECT 3.6500 1.4250 3.9100 1.5150 ;
      RECT 2.1500 1.4000 2.5800 1.4950 ;
      RECT 3.6500 0.8850 3.7400 1.4250 ;
      RECT 2.4900 1.0850 2.5800 1.4000 ;
      RECT 2.3850 0.9950 2.5800 1.0850 ;
      RECT 4.9600 1.9000 5.1500 1.9900 ;
      RECT 5.0550 0.6600 5.1500 1.9000 ;
      RECT 4.5050 0.5700 5.1500 0.6600 ;
      RECT 5.0300 0.4100 5.1500 0.5700 ;
      RECT 4.5050 0.6600 4.5950 1.2950 ;
      RECT 2.4900 0.4800 4.5950 0.5700 ;
      RECT 2.4900 0.5700 2.5800 0.8150 ;
      RECT 3.8300 0.5700 3.9200 1.3150 ;
      RECT 2.1800 0.8150 2.5800 0.9050 ;
      RECT 2.1800 0.9050 2.2700 1.2850 ;
  END
END DFFQ_X4M_A12TH

MACRO DFFRPQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8600 ;
        RECT 4.2750 0.3200 4.4450 0.8400 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 1.4100 3.9000 1.7100 ;
        RECT 3.8000 0.7750 3.9000 1.4100 ;
        RECT 3.7100 0.6750 3.9000 0.7750 ;
    END
    ANTENNADIFFAREA 0.151625 ;
  END QN

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7650 1.3900 ;
    END
    ANTENNAGATEAREA 0.0525 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.0750 1.5000 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.1600 1.4000 ;
    END
    ANTENNAGATEAREA 0.0192 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9850 4.5500 1.4050 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.2850 1.5200 0.4300 1.7100 ;
      RECT 0.2850 0.8600 0.3750 1.5200 ;
      RECT 0.2850 0.6500 0.4300 0.8600 ;
      RECT 0.5650 1.5750 0.8100 1.6650 ;
      RECT 0.7200 0.9400 0.8100 1.5750 ;
      RECT 0.7200 0.8500 1.3700 0.9400 ;
      RECT 1.2800 0.9400 1.3700 1.3950 ;
      RECT 0.7200 0.6700 0.8100 0.8500 ;
      RECT 0.9900 1.5700 2.0050 1.6600 ;
      RECT 1.9150 0.7500 2.0050 1.5700 ;
      RECT 1.5150 0.6600 2.0050 0.7500 ;
      RECT 0.9900 1.2400 1.0800 1.5700 ;
      RECT 3.1950 1.0600 3.2850 1.3300 ;
      RECT 2.6550 0.9900 3.2850 1.0600 ;
      RECT 2.0950 0.9700 3.2850 0.9900 ;
      RECT 2.0950 0.9900 2.1850 1.6950 ;
      RECT 2.0950 0.9000 2.7450 0.9700 ;
      RECT 2.5650 1.5350 3.4650 1.6250 ;
      RECT 2.5650 1.2200 2.6550 1.5350 ;
      RECT 3.3750 0.7700 3.4650 1.5350 ;
      RECT 3.0700 0.6800 3.4650 0.7700 ;
      RECT 0.5200 0.4800 4.1200 0.5700 ;
      RECT 4.0300 0.5700 4.1200 1.7100 ;
      RECT 0.5200 0.5700 0.6100 1.4550 ;
      RECT 0.6700 1.8300 4.7200 1.9200 ;
      RECT 4.6300 1.6100 4.7200 1.8300 ;
      RECT 4.6300 1.5200 4.7500 1.6100 ;
      RECT 4.6600 0.8700 4.7500 1.5200 ;
      RECT 4.6300 0.6800 4.7500 0.8700 ;
      RECT 2.3050 1.1100 2.3950 1.8300 ;
  END
END DFFRPQN_X0P5M_A12TH

MACRO DFFRPQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7600 ;
        RECT 1.1400 0.3200 1.3500 0.3900 ;
        RECT 1.8050 0.3200 2.0150 0.3900 ;
        RECT 2.9800 0.3200 3.1900 0.3900 ;
        RECT 3.5550 0.3200 3.7250 0.3700 ;
        RECT 4.3550 0.3200 4.4550 0.8700 ;
    END
  END VSS

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.1900 ;
        RECT 1.5000 0.8500 1.7500 0.9500 ;
    END
    ANTENNAGATEAREA 0.0687 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.0750 1.6900 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0300 0.1600 1.4550 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.9850 3.7500 1.2500 ;
        RECT 3.6500 1.2500 3.8450 1.3500 ;
        RECT 3.6500 0.8850 3.9500 0.9850 ;
        RECT 3.7450 1.3500 3.8450 1.7000 ;
        RECT 3.8500 0.7400 3.9500 0.8850 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3350 1.0000 4.5500 1.2100 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6600 0.4300 1.7500 ;
      RECT 0.7050 1.1000 1.5300 1.1900 ;
      RECT 0.5500 1.5850 0.7950 1.6750 ;
      RECT 0.7050 1.1900 0.7950 1.5850 ;
      RECT 0.7050 0.6900 0.7950 1.1000 ;
      RECT 1.7550 1.4250 1.8450 1.7200 ;
      RECT 0.9050 1.3350 1.9900 1.4250 ;
      RECT 1.9000 1.0350 1.9900 1.3350 ;
      RECT 1.9000 0.9450 2.3100 1.0350 ;
      RECT 1.9000 0.7600 1.9900 0.9450 ;
      RECT 1.4750 0.6700 1.9900 0.7600 ;
      RECT 1.9550 1.6200 2.5250 1.7100 ;
      RECT 2.4350 0.8550 2.5250 1.6200 ;
      RECT 2.4350 0.7650 3.2300 0.8550 ;
      RECT 3.1400 0.8550 3.2300 1.2900 ;
      RECT 2.4350 0.7600 2.5250 0.7650 ;
      RECT 2.1100 0.6700 2.5250 0.7600 ;
      RECT 2.8900 1.6100 3.5250 1.7000 ;
      RECT 2.8900 1.1200 2.9800 1.6100 ;
      RECT 3.4350 0.8650 3.5250 1.6100 ;
      RECT 3.3350 0.7750 3.5250 0.8650 ;
      RECT 4.0000 1.3000 4.1550 1.5100 ;
      RECT 4.0550 0.8400 4.1550 1.3000 ;
      RECT 4.0550 0.6700 4.1900 0.8400 ;
      RECT 4.0550 0.5800 4.1550 0.6700 ;
      RECT 0.5250 0.4900 4.1550 0.5800 ;
      RECT 0.5250 0.5800 0.6150 1.4750 ;
      RECT 0.7250 1.8300 4.7450 1.9200 ;
      RECT 4.6550 1.5400 4.7450 1.8300 ;
      RECT 4.6300 1.3300 4.7450 1.5400 ;
      RECT 4.6550 0.8400 4.7450 1.3300 ;
      RECT 4.6300 0.6500 4.7450 0.8400 ;
      RECT 1.9000 1.9200 2.1100 1.9900 ;
      RECT 2.6500 0.9800 2.7400 1.8300 ;
  END
END DFFRPQN_X1M_A12TH

MACRO DFFRPQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8300 ;
        RECT 3.7550 0.3200 3.9250 0.3700 ;
        RECT 4.2750 0.3200 4.4450 0.3700 ;
        RECT 4.7550 0.3200 4.8550 0.8700 ;
    END
  END VSS

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.1900 ;
        RECT 1.3200 0.8500 1.7500 0.9500 ;
    END
    ANTENNAGATEAREA 0.0957 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 0.0750 1.6500 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1600 1.4550 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.7350 4.1500 1.2500 ;
        RECT 3.9450 1.2500 4.1500 1.3500 ;
        RECT 3.9450 1.3500 4.0450 1.7000 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7350 1.0000 4.9500 1.2100 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3400 0.4900 0.4300 1.7550 ;
      RECT 0.7050 1.1000 1.4600 1.1900 ;
      RECT 0.5700 1.5850 0.7950 1.6750 ;
      RECT 0.7050 1.1900 0.7950 1.5850 ;
      RECT 0.7050 0.6900 0.7950 1.1000 ;
      RECT 1.7150 1.4250 1.8850 1.6400 ;
      RECT 0.9050 1.3350 1.9900 1.4250 ;
      RECT 1.9000 1.0050 1.9900 1.3350 ;
      RECT 1.9000 0.9150 2.5600 1.0050 ;
      RECT 1.9000 0.7600 1.9900 0.9150 ;
      RECT 1.4850 0.6700 1.9900 0.7600 ;
      RECT 1.9750 1.6200 2.7600 1.7100 ;
      RECT 1.9750 1.5400 2.1450 1.6200 ;
      RECT 2.6700 0.7900 2.7600 1.6200 ;
      RECT 2.1200 0.7000 3.4300 0.7900 ;
      RECT 3.3400 0.7900 3.4300 1.2900 ;
      RECT 3.0900 1.5550 3.7250 1.6450 ;
      RECT 3.0900 1.0700 3.1800 1.5550 ;
      RECT 3.6350 0.8150 3.7250 1.5550 ;
      RECT 3.5550 0.7250 3.7250 0.8150 ;
      RECT 4.4000 1.2750 4.5500 1.4850 ;
      RECT 4.4500 0.8600 4.5500 1.2750 ;
      RECT 4.4500 0.6500 4.5900 0.8600 ;
      RECT 4.4500 0.5800 4.5500 0.6500 ;
      RECT 0.5250 0.4900 4.5500 0.5800 ;
      RECT 0.5250 0.5800 0.6150 1.4750 ;
      RECT 0.7250 1.8300 5.1450 1.9200 ;
      RECT 5.0550 1.5400 5.1450 1.8300 ;
      RECT 5.0300 1.3300 5.1450 1.5400 ;
      RECT 5.0550 0.8600 5.1450 1.3300 ;
      RECT 5.0300 0.6500 5.1450 0.8600 ;
      RECT 2.8600 0.9100 2.9500 1.8300 ;
  END
END DFFRPQN_X2M_A12TH

MACRO DFFRPQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7300 ;
        RECT 3.7550 0.3200 3.9250 0.3700 ;
        RECT 4.2750 0.3200 4.4450 0.3700 ;
        RECT 5.1550 0.3200 5.2550 0.8650 ;
    END
  END VSS

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.1900 ;
        RECT 1.3200 0.8500 1.7500 0.9500 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.0750 1.7300 0.1750 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1600 1.4550 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.8900 4.5650 1.2400 ;
        RECT 3.9500 1.2400 4.5650 1.3400 ;
        RECT 3.9950 0.7900 4.7250 0.8900 ;
        RECT 3.9500 1.3400 4.0500 1.7000 ;
        RECT 4.4650 1.3400 4.5650 1.7000 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1350 1.0000 5.3500 1.2100 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.3400 0.4900 0.4300 1.9200 ;
      RECT 0.7050 1.1000 1.4600 1.1900 ;
      RECT 0.5700 1.5850 0.7950 1.6750 ;
      RECT 0.7050 1.1900 0.7950 1.5850 ;
      RECT 0.7050 0.7000 0.7950 1.1000 ;
      RECT 1.7100 1.4250 1.8800 1.6400 ;
      RECT 0.9050 1.3350 1.9900 1.4250 ;
      RECT 1.9000 1.0050 1.9900 1.3350 ;
      RECT 1.9000 0.9150 2.5600 1.0050 ;
      RECT 1.9000 0.7600 1.9900 0.9150 ;
      RECT 1.4850 0.6700 1.9900 0.7600 ;
      RECT 2.4100 1.6250 2.5000 1.7300 ;
      RECT 1.9700 1.5350 2.7600 1.6250 ;
      RECT 2.6700 0.7900 2.7600 1.5350 ;
      RECT 2.1200 0.7000 3.4300 0.7900 ;
      RECT 3.3400 0.7900 3.4300 1.0900 ;
      RECT 3.3400 1.0900 3.6250 1.1800 ;
      RECT 3.0900 1.5550 3.8250 1.6450 ;
      RECT 3.0900 1.0700 3.1800 1.5550 ;
      RECT 3.7350 0.8150 3.8250 1.5550 ;
      RECT 3.5400 0.7250 3.8250 0.8150 ;
      RECT 4.8000 1.2950 4.9500 1.5050 ;
      RECT 4.8500 0.8650 4.9500 1.2950 ;
      RECT 4.8500 0.6550 4.9900 0.8650 ;
      RECT 4.8500 0.5800 4.9500 0.6550 ;
      RECT 0.5250 0.4900 4.9500 0.5800 ;
      RECT 0.5250 0.5800 0.6150 1.4750 ;
      RECT 0.7250 1.8300 5.5450 1.9200 ;
      RECT 5.4550 1.5200 5.5450 1.8300 ;
      RECT 5.4300 1.3500 5.5450 1.5200 ;
      RECT 5.4550 0.8600 5.5450 1.3500 ;
      RECT 5.4250 0.6500 5.5450 0.8600 ;
      RECT 2.8600 0.9100 2.9500 1.8300 ;
  END
END DFFRPQN_X3M_A12TH

MACRO DFFRPQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8750 ;
        RECT 4.5100 0.3200 4.6100 0.8850 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8100 1.4500 4.0800 1.5500 ;
        RECT 3.9800 1.5500 4.0800 1.7100 ;
        RECT 3.9800 0.6700 4.0800 1.4500 ;
    END
    ANTENNADIFFAREA 0.131375 ;
  END Q

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6450 0.9800 1.7550 1.4000 ;
    END
    ANTENNAGATEAREA 0.0588 ;
  END R

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0800 1.5200 0.1700 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1600 1.4050 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 1.0050 4.7250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK
  OBS
    LAYER M1 ;
      RECT 0.2850 1.5200 0.4300 1.6900 ;
      RECT 0.2850 0.8400 0.3750 1.5200 ;
      RECT 0.2850 0.6700 0.4300 0.8400 ;
      RECT 0.5400 1.5750 0.8100 1.6650 ;
      RECT 0.7200 1.1300 0.8100 1.5750 ;
      RECT 0.7200 1.0400 1.4900 1.1300 ;
      RECT 1.4000 1.1300 1.4900 1.4300 ;
      RECT 0.7200 0.6700 0.8100 1.0400 ;
      RECT 0.9800 1.5700 1.9900 1.6600 ;
      RECT 1.9000 0.7500 1.9900 1.5700 ;
      RECT 1.5000 0.6600 1.9900 0.7500 ;
      RECT 0.9800 1.2400 1.0700 1.5700 ;
      RECT 3.1800 1.2000 3.3900 1.2900 ;
      RECT 3.1800 0.7850 3.2700 1.2000 ;
      RECT 2.1350 0.6950 3.2700 0.7850 ;
      RECT 2.1350 0.7850 2.2250 1.6900 ;
      RECT 3.5950 1.0550 3.8650 1.1450 ;
      RECT 2.6700 1.5500 3.6850 1.6400 ;
      RECT 3.5950 1.1450 3.6850 1.5500 ;
      RECT 2.6700 1.0100 2.7600 1.5500 ;
      RECT 3.5950 0.9300 3.6850 1.0550 ;
      RECT 3.3750 0.8400 3.6850 0.9300 ;
      RECT 3.3750 0.6900 3.4650 0.8400 ;
      RECT 0.5200 0.4800 4.3200 0.5700 ;
      RECT 4.2300 0.5700 4.3200 1.7100 ;
      RECT 0.4950 1.2850 0.6100 1.4550 ;
      RECT 0.5200 0.5700 0.6100 1.2850 ;
      RECT 0.6450 1.8300 4.9200 1.9200 ;
      RECT 4.8300 0.6800 4.9200 1.8300 ;
      RECT 2.4150 1.0750 2.5050 1.8300 ;
  END
END DFFRPQ_X0P5M_A12TH

MACRO DFFRPQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8800 ;
        RECT 4.5100 0.3200 4.6100 0.8850 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 1.0050 4.7250 1.1950 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9900 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END D

  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6450 0.9800 1.7550 1.4000 ;
    END
    ANTENNAGATEAREA 0.0669 ;
  END R

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8100 1.4500 4.0750 1.5500 ;
        RECT 3.9750 1.5500 4.0750 1.7100 ;
        RECT 3.9750 0.6700 4.0750 1.4500 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.0800 1.5700 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.6900 0.4300 1.7400 ;
      RECT 0.5400 1.5550 0.8100 1.6450 ;
      RECT 0.7200 1.1300 0.8100 1.5550 ;
      RECT 0.7200 1.0400 1.4950 1.1300 ;
      RECT 1.4050 1.1300 1.4950 1.4300 ;
      RECT 0.7200 0.6700 0.8100 1.0400 ;
      RECT 0.9750 1.5700 1.9900 1.6600 ;
      RECT 1.9000 0.7500 1.9900 1.5700 ;
      RECT 1.5000 0.6600 1.9900 0.7500 ;
      RECT 0.9750 1.2400 1.0650 1.5700 ;
      RECT 3.1800 1.2000 3.4550 1.2900 ;
      RECT 3.1800 0.7850 3.2700 1.2000 ;
      RECT 2.1350 0.6950 3.2700 0.7850 ;
      RECT 2.1350 0.7850 2.2250 1.6900 ;
      RECT 3.5950 1.0550 3.8650 1.1450 ;
      RECT 2.6700 1.5500 3.6850 1.6400 ;
      RECT 3.5950 1.1450 3.6850 1.5500 ;
      RECT 2.6700 1.0100 2.7600 1.5500 ;
      RECT 3.5950 0.9300 3.6850 1.0550 ;
      RECT 3.3750 0.8400 3.6850 0.9300 ;
      RECT 3.3750 0.7050 3.4650 0.8400 ;
      RECT 0.5200 0.4800 4.3200 0.5700 ;
      RECT 4.2300 0.5700 4.3200 1.7100 ;
      RECT 0.5200 0.5700 0.6100 1.4450 ;
      RECT 0.6450 1.8300 4.9200 1.9200 ;
      RECT 4.8300 0.6800 4.9200 1.8300 ;
      RECT 2.4150 1.0750 2.5050 1.8300 ;
  END
END DFFRPQ_X1M_A12TH

MACRO BUF_X4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.5950 0.3200 0.6950 0.7300 ;
        RECT 1.1150 0.3200 1.2150 0.7250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
        RECT 1.6300 1.4400 1.7200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 0.9500 1.3500 ;
        RECT 0.3350 1.3500 0.4350 1.7200 ;
        RECT 0.8550 1.3500 0.9500 1.7200 ;
        RECT 0.2500 0.9500 0.3500 1.2500 ;
        RECT 0.2500 0.8500 0.9500 0.9500 ;
        RECT 0.3350 0.5150 0.4350 0.8500 ;
        RECT 0.8500 0.5150 0.9500 0.8500 ;
    END
    ANTENNADIFFAREA 0.5958 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 1.0500 1.7050 1.1550 ;
    END
    ANTENNAGATEAREA 0.0918 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.3650 1.5300 1.4650 1.8300 ;
      RECT 1.0400 1.4400 1.4650 1.5300 ;
      RECT 1.0400 0.8300 1.5000 0.9200 ;
      RECT 1.4000 0.4900 1.5000 0.8300 ;
      RECT 1.0400 1.1500 1.1300 1.4400 ;
      RECT 0.4700 1.0500 1.1300 1.1500 ;
      RECT 1.0400 0.9200 1.1300 1.0500 ;
  END
END BUF_X4B_A12TH

MACRO BUF_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.9500 ;
        RECT 0.7200 0.3200 0.8100 0.6300 ;
        RECT 1.2400 0.3200 1.3300 0.6300 ;
        RECT 1.7600 0.3200 1.8500 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1074 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.7200 1.7700 0.8100 2.0800 ;
        RECT 1.2400 1.7700 1.3300 2.0800 ;
        RECT 1.7600 1.7700 1.8500 2.0800 ;
        RECT 0.1250 1.3700 0.2150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.2500 ;
        RECT 0.9750 1.2500 1.7500 1.3500 ;
        RECT 0.9800 0.8500 1.7500 0.9500 ;
        RECT 0.9800 1.3500 1.0700 1.7200 ;
        RECT 1.5000 1.3500 1.5900 1.7200 ;
        RECT 0.9800 0.4850 1.0700 0.8500 ;
        RECT 1.5000 0.4850 1.5900 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.4650 1.1500 ;
      RECT 0.3850 1.3700 0.4750 1.7200 ;
      RECT 0.3850 0.4850 0.4750 0.8300 ;
      RECT 0.3850 1.2800 0.7900 1.3700 ;
      RECT 0.7000 1.1500 0.7900 1.2800 ;
      RECT 0.7000 0.9200 0.7900 1.0600 ;
      RECT 0.3850 0.8300 0.7900 0.9200 ;
  END
END BUF_X4M_A12TH

MACRO BUF_X5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.7700 ;
        RECT 0.6750 0.3200 0.8450 0.7400 ;
        RECT 1.1950 0.3200 1.3650 0.7400 ;
        RECT 1.7150 0.3200 1.8850 0.7400 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.114 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9500 2.1500 1.2500 ;
        RECT 0.9750 1.2500 2.1500 1.3500 ;
        RECT 0.9750 0.8500 2.1500 0.9500 ;
        RECT 0.9750 1.3500 1.0650 1.7050 ;
        RECT 1.4950 1.3500 1.5850 1.7050 ;
        RECT 2.0150 1.3500 2.1500 1.7200 ;
        RECT 0.9750 0.4450 1.0650 0.8500 ;
        RECT 1.4950 0.4450 1.5850 0.8500 ;
        RECT 2.0150 0.4450 2.1500 0.8500 ;
    END
    ANTENNADIFFAREA 0.784875 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.7150 1.7700 0.8050 2.0800 ;
        RECT 1.2350 1.7700 1.3250 2.0800 ;
        RECT 1.7550 1.7700 1.8450 2.0800 ;
        RECT 0.1250 1.4950 0.2150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.8100 1.1500 ;
      RECT 0.3850 1.3700 0.4750 1.7200 ;
      RECT 0.3850 0.6650 0.4750 0.8300 ;
      RECT 0.3850 1.2800 0.7900 1.3700 ;
      RECT 0.7000 1.1500 0.7900 1.2800 ;
      RECT 0.7000 0.9200 0.7900 1.0600 ;
      RECT 0.3850 0.8300 0.7900 0.9200 ;
  END
END BUF_X5B_A12TH

MACRO BUF_X5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.8550 ;
        RECT 0.7150 0.3200 0.8050 0.6300 ;
        RECT 1.2350 0.3200 1.3250 0.6300 ;
        RECT 1.7550 0.3200 1.8450 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1332 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.7150 1.7700 0.8050 2.0800 ;
        RECT 1.2350 1.7700 1.3250 2.0800 ;
        RECT 1.7550 1.7700 1.8450 2.0800 ;
        RECT 0.1250 1.4800 0.2150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9500 2.1500 1.2500 ;
        RECT 0.9750 1.2500 2.1500 1.3500 ;
        RECT 0.9750 0.8500 2.1500 0.9500 ;
        RECT 0.9750 1.3500 1.0650 1.7200 ;
        RECT 1.4950 1.3500 1.5850 1.7200 ;
        RECT 2.0150 1.3500 2.1050 1.7200 ;
        RECT 0.9750 0.4850 1.0650 0.8500 ;
        RECT 1.4950 0.4850 1.5850 0.8500 ;
        RECT 2.0150 0.4850 2.1050 0.8500 ;
    END
    ANTENNADIFFAREA 0.934375 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.8050 1.1500 ;
      RECT 0.3850 1.3600 0.4750 1.7200 ;
      RECT 0.3850 0.4850 0.4750 0.8300 ;
      RECT 0.3850 1.2700 0.7900 1.3600 ;
      RECT 0.7000 1.1500 0.7900 1.2700 ;
      RECT 0.7000 0.9200 0.7900 1.0600 ;
      RECT 0.3850 0.8300 0.7900 0.9200 ;
  END
END BUF_X5M_A12TH

MACRO BUF_X6B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1200 0.3200 0.2100 0.9200 ;
        RECT 0.6350 0.3200 0.7350 0.7250 ;
        RECT 1.1350 0.3200 1.3050 0.7600 ;
        RECT 1.6550 0.3200 1.8250 0.7600 ;
        RECT 2.2150 0.3200 2.3050 0.8650 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1150 1.0500 0.5350 1.1500 ;
    END
    ANTENNAGATEAREA 0.1362 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.1750 1.7700 1.2650 2.0800 ;
        RECT 1.6950 1.7700 1.7850 2.0800 ;
        RECT 2.2150 1.7700 2.3050 2.0800 ;
        RECT 0.1200 1.6150 0.2100 2.0800 ;
        RECT 0.6400 1.6150 0.7300 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.2500 ;
        RECT 0.9150 1.2500 2.0450 1.3500 ;
        RECT 0.9150 0.8500 2.0450 0.9500 ;
        RECT 0.9150 1.3500 1.0050 1.7200 ;
        RECT 1.4350 1.3500 1.5250 1.7200 ;
        RECT 1.9550 1.3500 2.0450 1.7200 ;
        RECT 0.9150 0.4800 1.0050 0.8500 ;
        RECT 1.4350 0.4800 1.5250 0.8500 ;
        RECT 1.9550 0.4800 2.0450 0.8500 ;
    END
    ANTENNADIFFAREA 0.819 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.7300 1.1500 ;
      RECT 0.3800 1.3700 0.4700 1.7200 ;
      RECT 0.3800 0.5050 0.4700 0.8300 ;
      RECT 0.3800 1.2800 0.7900 1.3700 ;
      RECT 0.7000 1.1500 0.7900 1.2800 ;
      RECT 0.7000 0.9200 0.7900 1.0600 ;
      RECT 0.3800 0.8300 0.7900 0.9200 ;
  END
END BUF_X6B_A12TH

MACRO BUF_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1150 0.3200 0.2050 0.7600 ;
        RECT 0.6350 0.3200 0.7250 0.7400 ;
        RECT 1.1700 0.3200 1.2600 0.6200 ;
        RECT 1.6900 0.3200 1.7800 0.6200 ;
        RECT 2.2100 0.3200 2.3000 0.6200 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1100 1.0500 0.5300 1.1500 ;
    END
    ANTENNAGATEAREA 0.1596 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.1700 1.7700 1.2600 2.0800 ;
        RECT 1.6900 1.7700 1.7800 2.0800 ;
        RECT 2.2100 1.7700 2.3000 2.0800 ;
        RECT 0.1150 1.6050 0.2050 2.0800 ;
        RECT 0.6500 1.6050 0.7400 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9500 2.1500 1.2500 ;
        RECT 0.9100 1.2500 2.1500 1.3500 ;
        RECT 0.9100 0.8500 2.1500 0.9500 ;
        RECT 0.9100 1.3500 1.0000 1.7200 ;
        RECT 1.4300 1.3500 1.5200 1.7200 ;
        RECT 1.9500 1.3500 2.0400 1.7200 ;
        RECT 0.9100 0.4850 1.0000 0.8500 ;
        RECT 1.4300 0.4850 1.5200 0.8500 ;
        RECT 1.9500 0.4850 2.0400 0.8500 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0600 1.8500 1.1500 ;
      RECT 0.3750 1.3700 0.4650 1.7200 ;
      RECT 0.3750 0.4850 0.4650 0.8300 ;
      RECT 0.3750 1.2800 0.7900 1.3700 ;
      RECT 0.7000 1.1500 0.7900 1.2800 ;
      RECT 0.7000 0.9200 0.7900 1.0600 ;
      RECT 0.3750 0.8300 0.7900 0.9200 ;
  END
END BUF_X6M_A12TH

MACRO BUF_X7P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.7400 ;
        RECT 0.8650 0.3200 1.0350 0.7400 ;
        RECT 1.4350 0.3200 1.5350 0.7100 ;
        RECT 1.9550 0.3200 2.0550 0.7100 ;
        RECT 2.4750 0.3200 2.5750 0.7100 ;
        RECT 3.0000 0.3200 3.0900 0.9150 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 1.4400 1.7200 1.5300 2.0800 ;
        RECT 1.9600 1.7200 2.0500 2.0800 ;
        RECT 2.4800 1.7200 2.5700 2.0800 ;
        RECT 3.0000 1.7200 3.0900 2.0800 ;
        RECT 0.9050 1.5250 0.9950 2.0800 ;
        RECT 0.3850 1.5050 0.4750 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1737 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6450 0.9550 2.7550 1.2450 ;
        RECT 1.1800 1.2450 2.8300 1.3550 ;
        RECT 1.1800 0.8450 2.8300 0.9550 ;
        RECT 1.1800 1.3550 1.2700 1.7250 ;
        RECT 1.7000 1.3550 1.7900 1.7250 ;
        RECT 2.2200 1.3550 2.3100 1.7250 ;
        RECT 2.7400 1.3550 2.8300 1.7250 ;
        RECT 1.1800 0.4850 1.2700 0.8450 ;
        RECT 1.7000 0.4850 1.7900 0.8450 ;
        RECT 2.2200 0.4850 2.3100 0.8450 ;
        RECT 2.7400 0.4850 2.8300 0.8450 ;
    END
    ANTENNADIFFAREA 1.028 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.9200 1.0600 2.4150 1.1500 ;
      RECT 0.1250 1.3700 0.2150 1.7200 ;
      RECT 0.1250 0.7050 0.2150 0.8300 ;
      RECT 0.6450 1.3700 0.7350 1.7200 ;
      RECT 0.6450 0.7050 0.7350 0.8300 ;
      RECT 0.1250 1.2800 1.0100 1.3700 ;
      RECT 0.9200 1.1500 1.0100 1.2800 ;
      RECT 0.9200 0.9200 1.0100 1.0600 ;
      RECT 0.1250 0.8300 1.0100 0.9200 ;
  END
END BUF_X7P5B_A12TH

MACRO BUF_X7P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.1400 0.3200 0.2400 0.6900 ;
        RECT 0.6600 0.3200 0.7600 0.7250 ;
        RECT 1.2050 0.3200 1.3050 0.7300 ;
        RECT 1.7250 0.3200 1.8250 0.7300 ;
        RECT 2.2450 0.3200 2.3450 0.7300 ;
        RECT 2.7650 0.3200 2.8650 0.7300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 0.9600 2.7600 1.4400 ;
        RECT 0.9350 1.4400 2.7600 1.5600 ;
        RECT 0.9350 0.8400 2.7600 0.9600 ;
        RECT 0.9350 1.5600 1.0550 1.8950 ;
        RECT 1.4550 1.5600 1.5750 1.8400 ;
        RECT 1.9750 1.5600 2.0950 1.8400 ;
        RECT 2.4950 1.5600 2.6150 1.8400 ;
        RECT 1.4550 0.5300 1.5750 0.8400 ;
        RECT 1.9750 0.5300 2.0950 0.8400 ;
        RECT 2.4950 0.5300 2.6150 0.8400 ;
        RECT 0.9350 0.5250 1.0550 0.8400 ;
    END
    ANTENNADIFFAREA 1.224 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.0500 0.6300 1.1500 ;
    END
    ANTENNAGATEAREA 0.195 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.1400 1.7550 0.2400 2.0800 ;
        RECT 0.6600 1.7100 0.7600 2.0800 ;
        RECT 1.2050 1.7100 1.3050 2.0800 ;
        RECT 1.7250 1.7100 1.8250 2.0800 ;
        RECT 2.2450 1.7100 2.3450 2.0800 ;
        RECT 2.7650 1.7100 2.8650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7400 1.0900 1.7450 1.1800 ;
      RECT 0.4050 1.5500 0.4950 1.9150 ;
      RECT 0.4050 0.5200 0.4950 0.8400 ;
      RECT 0.4050 1.4600 0.8300 1.5500 ;
      RECT 0.7400 1.1800 0.8300 1.4600 ;
      RECT 0.7400 0.9300 0.8300 1.0900 ;
      RECT 0.4050 0.8400 0.8300 0.9300 ;
  END
END BUF_X7P5M_A12TH

MACRO BUF_X9B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.2800 0.3200 0.3700 0.7750 ;
        RECT 0.8000 0.3200 0.8900 0.7400 ;
        RECT 1.3900 0.3200 1.4900 0.6700 ;
        RECT 1.9100 0.3200 2.0100 0.6700 ;
        RECT 2.4300 0.3200 2.5300 0.6700 ;
        RECT 2.9500 0.3200 3.0500 0.6700 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
        RECT 1.9150 1.7700 2.0050 2.0800 ;
        RECT 2.4350 1.7700 2.5250 2.0800 ;
        RECT 2.9550 1.7700 3.0450 2.0800 ;
        RECT 0.3550 1.6400 0.4450 2.0800 ;
        RECT 0.8750 1.6400 0.9650 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1350 1.2350 3.3050 1.3650 ;
        RECT 1.1350 1.3650 1.2250 1.7200 ;
        RECT 1.6550 1.3650 1.7450 1.7200 ;
        RECT 2.1750 1.3650 2.2650 1.7200 ;
        RECT 2.6950 1.3650 2.7850 1.7200 ;
        RECT 3.2150 1.3650 3.3050 1.7200 ;
        RECT 3.0350 0.9650 3.1650 1.2350 ;
        RECT 1.1350 0.8350 3.3050 0.9650 ;
        RECT 1.1350 0.4850 1.2250 0.8350 ;
        RECT 1.6550 0.4850 1.7450 0.8350 ;
        RECT 2.1750 0.4850 2.2650 0.8350 ;
        RECT 2.6950 0.4850 2.7850 0.8350 ;
        RECT 3.2150 0.4850 3.3050 0.8350 ;
    END
    ANTENNADIFFAREA 1.330875 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 0.7300 1.1500 ;
    END
    ANTENNAGATEAREA 0.2052 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.9000 1.0550 2.7750 1.1450 ;
      RECT 0.6150 1.3700 0.7050 1.7200 ;
      RECT 0.5400 0.4850 0.6300 0.8300 ;
      RECT 0.0950 1.2800 0.9900 1.3700 ;
      RECT 0.9000 1.1450 0.9900 1.2800 ;
      RECT 0.9000 0.9200 0.9900 1.0550 ;
      RECT 0.5400 0.8300 0.9900 0.9200 ;
      RECT 0.0950 1.3700 0.1850 1.7200 ;
  END
END BUF_X9B_A12TH

MACRO BUF_X9M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7350 ;
        RECT 0.8750 0.3200 0.9650 0.7350 ;
        RECT 1.3950 0.3200 1.4850 0.6300 ;
        RECT 1.9150 0.3200 2.0050 0.6300 ;
        RECT 2.4350 0.3200 2.5250 0.6300 ;
        RECT 2.9550 0.3200 3.0450 0.6300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1350 1.2350 3.3050 1.3650 ;
        RECT 1.1350 1.3650 1.2250 1.7200 ;
        RECT 1.6550 1.3650 1.7450 1.7200 ;
        RECT 2.1750 1.3650 2.2650 1.7200 ;
        RECT 2.6950 1.3650 2.7850 1.7200 ;
        RECT 3.2150 1.3650 3.3050 1.7200 ;
        RECT 3.0350 0.9650 3.1650 1.2350 ;
        RECT 1.1350 0.8350 3.3050 0.9650 ;
        RECT 1.1350 0.5050 1.2250 0.8350 ;
        RECT 1.6550 0.5050 1.7450 0.8350 ;
        RECT 2.1750 0.5050 2.2650 0.8350 ;
        RECT 2.6950 0.5050 2.7850 0.8350 ;
        RECT 3.2150 0.5050 3.3050 0.8350 ;
    END
    ANTENNADIFFAREA 1.584375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 1.0500 0.7550 1.1500 ;
    END
    ANTENNAGATEAREA 0.2412 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
        RECT 1.9150 1.7700 2.0050 2.0800 ;
        RECT 2.4350 1.7700 2.5250 2.0800 ;
        RECT 2.9550 1.7700 3.0450 2.0800 ;
        RECT 0.3550 1.6100 0.4450 2.0800 ;
        RECT 0.8750 1.6100 0.9650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.9000 1.0550 2.7500 1.1450 ;
      RECT 0.0950 1.2800 0.9900 1.3700 ;
      RECT 0.9000 1.1450 0.9900 1.2800 ;
      RECT 0.9000 0.9200 0.9900 1.0550 ;
      RECT 0.0950 0.8300 0.9900 0.9200 ;
      RECT 0.0950 1.3700 0.1850 1.7200 ;
      RECT 0.0950 0.4850 0.1850 0.8300 ;
      RECT 0.6150 1.3700 0.7050 1.7200 ;
      RECT 0.6150 0.4850 0.7050 0.8300 ;
  END
END BUF_X9M_A12TH

MACRO CGENCIN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 3.8250 1.7450 3.9250 2.0800 ;
    END
  END VDD

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.8100 3.7850 1.1900 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END CIN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9150 1.0500 1.5100 1.1500 ;
        RECT 1.4100 1.1500 1.5100 1.2850 ;
        RECT 1.4100 0.9600 1.5100 1.0500 ;
        RECT 1.4100 1.2850 1.6400 1.3800 ;
        RECT 1.4100 0.8600 2.3150 0.9600 ;
        RECT 2.2250 0.9600 2.3150 1.0850 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 1.2500 1.1900 1.3500 ;
        RECT 0.6300 1.0200 0.7400 1.2500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2400 0.7100 3.3800 1.3800 ;
        RECT 3.1250 0.6200 3.3800 0.7100 ;
        RECT 3.1250 0.4850 3.2150 0.6200 ;
    END
    ANTENNADIFFAREA 0.2321 ;
  END CO

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3050 0.3200 0.6750 0.3750 ;
        RECT 2.3400 0.3200 2.5500 0.3900 ;
        RECT 3.6800 0.3200 3.7850 0.7050 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.8800 1.6500 3.0450 1.7400 ;
      RECT 0.4450 0.9300 0.5350 1.4700 ;
      RECT 0.4450 0.8400 1.2700 0.9300 ;
      RECT 1.8800 1.5600 1.9700 1.6500 ;
      RECT 0.4450 1.4700 1.9700 1.5600 ;
      RECT 1.3200 1.8800 3.5900 1.9200 ;
      RECT 3.3250 1.9200 3.5900 1.9700 ;
      RECT 1.3200 1.8300 3.4400 1.8800 ;
      RECT 3.3500 1.5600 3.4400 1.8300 ;
      RECT 2.9450 1.4700 3.4400 1.5600 ;
      RECT 2.9450 0.5700 3.0350 1.4700 ;
      RECT 1.5800 0.4800 3.0350 0.5700 ;
      RECT 1.3200 1.9200 1.4900 1.9400 ;
      RECT 1.5800 0.4600 1.7700 0.4800 ;
      RECT 3.5650 1.3700 3.6550 1.7300 ;
      RECT 3.4700 1.2800 3.6550 1.3700 ;
      RECT 3.4700 0.5300 3.5600 1.2800 ;
      RECT 3.3300 0.4400 3.5600 0.5300 ;
      RECT 0.0450 0.4800 1.4900 0.5700 ;
      RECT 1.3000 0.4600 1.4900 0.4800 ;
      RECT 0.0450 1.3900 0.1700 1.8300 ;
      RECT 0.0450 0.7050 0.1350 1.3900 ;
      RECT 0.0450 0.5700 0.1700 0.7050 ;
      RECT 1.0600 1.9200 1.2300 1.9400 ;
      RECT 0.0450 1.8300 1.2300 1.9200 ;
      RECT 0.2650 1.6500 1.7700 1.7400 ;
      RECT 0.2650 0.6600 2.0100 0.7500 ;
      RECT 1.8350 0.7500 2.0100 0.7700 ;
      RECT 0.2650 1.1550 0.3550 1.6500 ;
      RECT 0.2300 0.9050 0.3550 1.1550 ;
      RECT 0.2650 0.7500 0.3550 0.9050 ;
      RECT 2.1400 1.3300 2.2300 1.5250 ;
      RECT 1.9650 1.2400 2.5650 1.3300 ;
      RECT 2.4750 0.7500 2.5650 1.2400 ;
      RECT 2.1000 0.6600 2.5650 0.7500 ;
      RECT 2.1000 0.7500 2.2750 0.7700 ;
      RECT 1.9650 1.1500 2.0550 1.2400 ;
      RECT 1.7150 1.0500 2.0550 1.1500 ;
      RECT 2.7550 0.7700 2.8550 1.4950 ;
      RECT 2.6550 0.6600 2.8550 0.7700 ;
  END
END CGENCIN_X1M_A12TH

MACRO CGENCIN_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 5.0600 2.0200 5.1700 2.0800 ;
        RECT 5.5950 2.0150 5.7050 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 1.0450 0.7550 1.2500 ;
        RECT 0.6200 1.2500 1.1900 1.3500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2150 0.8750 5.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.1212 ;
  END CIN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9350 1.0500 1.6200 1.1500 ;
        RECT 1.5200 1.1500 1.6200 1.2500 ;
        RECT 1.5200 0.9500 1.6200 1.0500 ;
        RECT 1.5200 1.2500 1.8250 1.3500 ;
        RECT 1.5200 0.8400 1.7500 0.9500 ;
        RECT 1.7250 1.3500 1.8250 1.4600 ;
        RECT 1.7250 1.4600 2.2350 1.5600 ;
        RECT 2.1350 1.2000 2.2350 1.4600 ;
        RECT 2.1350 1.1100 2.6750 1.2000 ;
    END
    ANTENNAGATEAREA 0.2412 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.2900 0.3200 0.7100 0.3700 ;
        RECT 2.4450 0.3200 2.5450 0.5400 ;
        RECT 2.9650 0.3200 3.0650 0.5400 ;
        RECT 3.5050 0.3200 3.6050 0.5400 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7200 1.6500 5.0100 1.7500 ;
        RECT 4.9100 1.7500 5.0100 1.8200 ;
        RECT 4.9100 1.8200 5.7500 1.9200 ;
        RECT 5.6500 0.5800 5.7500 1.8200 ;
        RECT 3.7200 0.4800 5.7500 0.5800 ;
    END
    ANTENNADIFFAREA 0.364 ;
  END CO
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5400 0.5700 ;
      RECT 1.3250 0.4600 1.5400 0.4800 ;
      RECT 0.0450 1.3900 0.1700 1.8300 ;
      RECT 0.0450 0.6900 0.1350 1.3900 ;
      RECT 0.0450 0.5700 0.1700 0.6900 ;
      RECT 0.0450 1.8300 1.2500 1.9200 ;
      RECT 0.2600 0.6600 2.0100 0.7500 ;
      RECT 1.9200 0.7500 2.0100 1.1300 ;
      RECT 1.9200 1.1300 2.0300 1.3700 ;
      RECT 0.2600 1.6400 0.7300 1.7300 ;
      RECT 0.2600 1.1550 0.3500 1.6400 ;
      RECT 0.2300 0.9050 0.3500 1.1550 ;
      RECT 0.2600 0.7500 0.3500 0.9050 ;
      RECT 2.6400 1.4700 3.0650 1.5600 ;
      RECT 2.9750 1.0300 3.0650 1.4700 ;
      RECT 2.9750 0.9300 3.4950 1.0300 ;
      RECT 2.9750 0.8400 3.0650 0.9300 ;
      RECT 2.3100 0.7500 3.0650 0.8400 ;
      RECT 2.3100 0.7300 2.8100 0.7500 ;
      RECT 2.7000 0.4500 2.8100 0.7300 ;
      RECT 3.5750 1.9200 3.9950 1.9600 ;
      RECT 1.3450 1.8700 3.9950 1.9200 ;
      RECT 1.3450 1.8300 3.6650 1.8700 ;
      RECT 0.4400 0.9300 0.5300 1.4600 ;
      RECT 1.3450 1.7100 1.4350 1.8300 ;
      RECT 0.8500 1.6200 1.4350 1.7100 ;
      RECT 0.8500 1.5500 0.9400 1.6200 ;
      RECT 0.4400 1.4600 0.9400 1.5500 ;
      RECT 0.4400 0.8400 1.3000 0.9300 ;
      RECT 3.2150 1.2900 4.1950 1.3800 ;
      RECT 3.5850 1.2700 4.1950 1.2900 ;
      RECT 3.2400 0.6700 4.2050 0.7600 ;
      RECT 3.5850 0.7600 3.6850 1.2700 ;
      RECT 3.2150 1.3800 3.3750 1.4850 ;
      RECT 3.2400 0.4650 3.3400 0.6700 ;
      RECT 3.4900 1.4700 4.3850 1.5600 ;
      RECT 4.2950 1.2550 4.3850 1.4700 ;
      RECT 4.2950 1.1650 4.8750 1.2550 ;
      RECT 4.2950 0.9650 4.3850 1.1650 ;
      RECT 3.8500 0.8750 4.3850 0.9650 ;
      RECT 1.5450 1.6500 3.5800 1.7400 ;
      RECT 3.4900 1.5600 3.5800 1.6500 ;
      RECT 2.1100 0.6200 2.2000 0.9300 ;
      RECT 2.1100 0.5700 2.3050 0.6200 ;
      RECT 1.6300 0.4800 2.3050 0.5700 ;
      RECT 1.5450 1.5300 1.6350 1.6500 ;
      RECT 1.3200 1.4400 1.6350 1.5300 ;
      RECT 1.6300 0.4600 1.8400 0.4800 ;
      RECT 2.3550 1.3800 2.4450 1.6500 ;
      RECT 2.3550 1.2900 2.8750 1.3800 ;
      RECT 2.7850 1.0200 2.8750 1.2900 ;
      RECT 2.1100 0.9300 2.8750 1.0200 ;
      RECT 5.3100 1.5300 5.4700 1.7300 ;
      RECT 4.4850 1.4300 5.5600 1.5300 ;
      RECT 5.4700 0.7600 5.5600 1.4300 ;
      RECT 4.4850 0.6700 5.5600 0.7600 ;
  END
END CGENCIN_X1P4M_A12TH

MACRO CGENCIN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 5.0400 1.9650 5.1500 2.0800 ;
        RECT 5.5750 1.9600 5.6850 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 1.2500 1.1900 1.3500 ;
        RECT 0.6200 1.0450 0.7550 1.2500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2150 0.8750 5.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.168 ;
  END CIN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9350 1.0500 1.6200 1.1500 ;
        RECT 1.5200 1.1500 1.6200 1.2500 ;
        RECT 1.5200 0.9500 1.6200 1.0500 ;
        RECT 1.5200 1.2500 1.8250 1.3500 ;
        RECT 1.5200 0.8400 1.7500 0.9500 ;
        RECT 1.7250 1.3500 1.8250 1.4600 ;
        RECT 1.7250 1.4600 2.2350 1.5600 ;
        RECT 2.1350 1.2000 2.2350 1.4600 ;
        RECT 2.1350 1.1100 2.6750 1.2000 ;
    END
    ANTENNAGATEAREA 0.2844 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.2900 0.3200 0.7000 0.3700 ;
        RECT 2.4450 0.3200 2.5450 0.6400 ;
        RECT 2.9650 0.3200 3.0650 0.6400 ;
        RECT 3.4650 0.3200 3.6050 0.5450 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7000 1.6500 4.8900 1.7500 ;
        RECT 4.7900 1.7500 4.8900 1.7600 ;
        RECT 4.7900 1.7600 5.7500 1.8600 ;
        RECT 5.6500 0.5800 5.7500 1.7600 ;
        RECT 3.7000 0.4800 5.7500 0.5800 ;
        RECT 3.7000 0.4700 3.9150 0.4800 ;
    END
    ANTENNADIFFAREA 0.52805 ;
  END CO
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5400 0.5700 ;
      RECT 1.3250 0.4600 1.5400 0.4800 ;
      RECT 0.0450 1.3900 0.1700 1.8300 ;
      RECT 0.0450 0.6900 0.1350 1.3900 ;
      RECT 0.0450 0.5700 0.1700 0.6900 ;
      RECT 0.0450 1.8300 1.2500 1.9200 ;
      RECT 0.2600 0.6600 2.0100 0.7500 ;
      RECT 1.9200 0.7500 2.0100 1.1300 ;
      RECT 1.9200 1.1300 2.0300 1.3700 ;
      RECT 0.2600 1.6400 0.7300 1.7300 ;
      RECT 0.2600 1.1550 0.3500 1.6400 ;
      RECT 0.2300 0.9050 0.3500 1.1550 ;
      RECT 0.2600 0.7500 0.3500 0.9050 ;
      RECT 2.9750 0.9300 3.4750 1.0300 ;
      RECT 2.3100 0.7300 2.8100 0.7500 ;
      RECT 2.7000 0.4500 2.8100 0.7300 ;
      RECT 2.6400 1.4700 3.0650 1.5600 ;
      RECT 2.9750 1.0300 3.0650 1.4700 ;
      RECT 2.9750 0.8400 3.0650 0.9300 ;
      RECT 2.3100 0.7500 3.0650 0.8400 ;
      RECT 3.5550 1.9200 3.9750 1.9600 ;
      RECT 1.3450 1.8700 3.9750 1.9200 ;
      RECT 1.3450 1.8300 3.6450 1.8700 ;
      RECT 0.4400 0.9300 0.5300 1.4600 ;
      RECT 1.3450 1.7100 1.4350 1.8300 ;
      RECT 0.8500 1.6200 1.4350 1.7100 ;
      RECT 0.8500 1.5500 0.9400 1.6200 ;
      RECT 0.4400 1.4600 0.9400 1.5500 ;
      RECT 0.4400 0.8400 1.3000 0.9300 ;
      RECT 3.1950 1.2900 4.1750 1.3800 ;
      RECT 3.5650 1.2700 4.1750 1.2900 ;
      RECT 3.2200 0.6700 4.1850 0.7600 ;
      RECT 3.5650 0.7600 3.6650 1.2700 ;
      RECT 3.1950 1.3800 3.3550 1.4850 ;
      RECT 3.2200 0.4650 3.3200 0.6700 ;
      RECT 3.4700 1.4700 4.3650 1.5600 ;
      RECT 4.2750 1.2550 4.3650 1.4700 ;
      RECT 4.2750 1.1650 4.8550 1.2550 ;
      RECT 4.2750 0.9650 4.3650 1.1650 ;
      RECT 3.8150 0.8750 4.3650 0.9650 ;
      RECT 1.5450 1.6500 3.5600 1.7400 ;
      RECT 3.4700 1.5600 3.5600 1.6500 ;
      RECT 2.1100 0.6200 2.2000 0.9300 ;
      RECT 2.1100 0.5700 2.3050 0.6200 ;
      RECT 1.6300 0.4800 2.3050 0.5700 ;
      RECT 1.5450 1.5300 1.6350 1.6500 ;
      RECT 1.3200 1.4400 1.6350 1.5300 ;
      RECT 1.6300 0.4600 1.8400 0.4800 ;
      RECT 2.3550 1.3800 2.4450 1.6500 ;
      RECT 2.3550 1.2900 2.8750 1.3800 ;
      RECT 2.7850 1.0200 2.8750 1.2900 ;
      RECT 2.1100 0.9300 2.8750 1.0200 ;
      RECT 5.2900 1.5250 5.4500 1.6700 ;
      RECT 4.4650 1.4250 5.4500 1.5250 ;
      RECT 5.2900 1.3850 5.4500 1.4250 ;
      RECT 5.2900 1.2850 5.5600 1.3850 ;
      RECT 5.4700 0.7600 5.5600 1.2850 ;
      RECT 4.4650 0.6700 5.5600 0.7600 ;
  END
END CGENCIN_X2M_A12TH

MACRO CGENCON_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 3.4250 1.7450 3.5250 2.0800 ;
    END
  END VDD

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.8100 3.3850 1.1900 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END CI

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9150 1.0500 1.5100 1.1500 ;
        RECT 1.4100 1.1500 1.5100 1.2850 ;
        RECT 1.4100 0.9500 1.5100 1.0500 ;
        RECT 1.4100 1.2850 1.6500 1.3800 ;
        RECT 1.4100 0.8500 2.2650 0.9500 ;
        RECT 2.0750 0.8400 2.2650 0.8500 ;
    END
    ANTENNAGATEAREA 0.2046 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.3050 0.3200 0.6750 0.3750 ;
        RECT 3.2800 0.3200 3.3850 0.7050 ;
    END
  END VSS

  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8400 0.7100 2.9800 1.3800 ;
        RECT 2.7250 0.6200 2.9800 0.7100 ;
        RECT 2.7250 0.4850 2.8150 0.6200 ;
    END
    ANTENNADIFFAREA 0.2321 ;
  END CON

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 1.2500 1.1900 1.3500 ;
        RECT 0.6300 1.0200 0.7400 1.2500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.4900 0.5700 ;
      RECT 1.3000 0.4600 1.4900 0.4800 ;
      RECT 0.0450 1.3900 0.1700 1.8300 ;
      RECT 0.0450 0.7950 0.1350 1.3900 ;
      RECT 0.0450 0.5700 0.1700 0.7950 ;
      RECT 1.0600 1.9200 1.2300 1.9400 ;
      RECT 0.0450 1.8300 1.2300 1.9200 ;
      RECT 0.2650 1.6500 1.7550 1.7400 ;
      RECT 0.2650 0.6600 2.0300 0.7500 ;
      RECT 0.2650 1.1550 0.3550 1.6500 ;
      RECT 0.2300 0.9050 0.3550 1.1550 ;
      RECT 0.2650 0.7500 0.3550 0.9050 ;
      RECT 2.3550 1.1500 2.4550 1.4950 ;
      RECT 1.7150 1.0500 2.4550 1.1500 ;
      RECT 2.3550 0.6800 2.4550 1.0500 ;
      RECT 1.8800 1.6500 2.6450 1.7400 ;
      RECT 0.4450 0.9300 0.5350 1.4700 ;
      RECT 0.4450 0.8400 1.2700 0.9300 ;
      RECT 1.8800 1.5600 1.9700 1.6500 ;
      RECT 0.4450 1.4700 1.9700 1.5600 ;
      RECT 1.3200 1.8800 3.1900 1.9200 ;
      RECT 2.9250 1.9200 3.1900 1.9700 ;
      RECT 1.3200 1.8300 3.0400 1.8800 ;
      RECT 2.9500 1.5600 3.0400 1.8300 ;
      RECT 2.5450 1.4700 3.0400 1.5600 ;
      RECT 2.5450 0.5700 2.6350 1.4700 ;
      RECT 1.5800 0.4800 2.6350 0.5700 ;
      RECT 1.3200 1.9200 1.4900 1.9400 ;
      RECT 1.5800 0.4600 1.7700 0.4800 ;
      RECT 3.1650 1.3700 3.2550 1.7200 ;
      RECT 3.0700 1.2800 3.2550 1.3700 ;
      RECT 3.0700 0.5300 3.1600 1.2800 ;
      RECT 2.9300 0.4400 3.1600 0.5300 ;
  END
END CGENCON_X1M_A12TH

MACRO CGENCON_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 4.4750 1.9650 4.5850 2.0800 ;
        RECT 5.0100 1.9600 5.1200 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 1.0450 0.7550 1.2500 ;
        RECT 0.6200 1.2500 1.1700 1.3500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6150 0.8750 4.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.1212 ;
  END CI

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9150 1.0500 1.6000 1.1500 ;
        RECT 1.5000 1.1500 1.6000 1.2500 ;
        RECT 1.5000 0.9500 1.6000 1.0500 ;
        RECT 1.5000 1.2500 1.8050 1.3500 ;
        RECT 1.5000 0.8400 1.7300 0.9500 ;
        RECT 1.7050 1.3500 1.8050 1.4600 ;
        RECT 1.7050 1.4600 2.2150 1.5600 ;
        RECT 2.1150 1.2200 2.2150 1.4600 ;
        RECT 2.1150 1.1100 2.3800 1.2200 ;
    END
    ANTENNAGATEAREA 0.2412 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.2750 0.3200 0.6950 0.3700 ;
        RECT 2.4050 0.3200 2.5050 0.5400 ;
        RECT 2.9250 0.3200 3.0250 0.5400 ;
    END
  END VSS

  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1200 1.6500 4.4050 1.7500 ;
        RECT 4.3050 1.7500 4.4050 1.7600 ;
        RECT 4.3050 1.7600 5.1500 1.8600 ;
        RECT 5.0500 0.5800 5.1500 1.7600 ;
        RECT 3.1200 0.4800 5.1500 0.5800 ;
        RECT 3.1200 0.4700 3.3350 0.4800 ;
    END
    ANTENNADIFFAREA 0.350925 ;
  END CON
  OBS
    LAYER M1 ;
      RECT 0.2600 0.6600 1.9900 0.7500 ;
      RECT 1.9000 0.7500 1.9900 1.1300 ;
      RECT 1.9000 1.1300 2.0100 1.3700 ;
      RECT 0.2600 1.6200 0.7300 1.7300 ;
      RECT 0.2600 1.1550 0.3500 1.6200 ;
      RECT 0.2300 0.9050 0.3500 1.1550 ;
      RECT 0.2600 0.7500 0.3500 0.9050 ;
      RECT 2.9750 1.9200 3.3950 1.9600 ;
      RECT 1.3250 1.8700 3.3950 1.9200 ;
      RECT 1.3250 1.8300 3.0650 1.8700 ;
      RECT 1.3250 1.7100 1.4150 1.8300 ;
      RECT 0.8300 1.6200 1.4150 1.7100 ;
      RECT 0.8300 1.5300 0.9400 1.6200 ;
      RECT 0.4400 1.4400 0.9400 1.5300 ;
      RECT 0.4400 0.8400 1.2800 0.9300 ;
      RECT 0.4400 0.9300 0.5300 1.4400 ;
      RECT 2.6600 1.2900 3.5950 1.3800 ;
      RECT 3.3400 1.2700 3.5950 1.2900 ;
      RECT 2.2900 0.7300 3.6050 0.7600 ;
      RECT 2.6600 0.6700 3.6050 0.7300 ;
      RECT 2.6600 1.3800 2.7700 1.5600 ;
      RECT 2.6600 0.8400 2.7500 1.2900 ;
      RECT 2.2900 0.7600 2.7500 0.8400 ;
      RECT 2.6600 0.4500 2.7700 0.6700 ;
      RECT 2.9100 1.4700 3.7850 1.5600 ;
      RECT 3.6950 1.2550 3.7850 1.4700 ;
      RECT 3.6950 1.1650 4.2750 1.2550 ;
      RECT 3.6950 0.9650 3.7850 1.1650 ;
      RECT 3.2500 0.8750 3.7850 0.9650 ;
      RECT 1.5250 1.6500 3.0000 1.7400 ;
      RECT 2.9100 1.5600 3.0000 1.6500 ;
      RECT 2.0900 0.6200 2.1800 0.9300 ;
      RECT 2.0900 0.5700 2.2850 0.6200 ;
      RECT 1.6100 0.4800 2.2850 0.5700 ;
      RECT 1.5250 1.5300 1.6150 1.6500 ;
      RECT 1.3000 1.4400 1.6150 1.5300 ;
      RECT 1.6100 0.4600 1.8200 0.4800 ;
      RECT 2.4700 1.0200 2.5600 1.6500 ;
      RECT 2.0900 0.9300 2.5600 1.0200 ;
      RECT 4.7250 1.5400 4.8850 1.6700 ;
      RECT 3.9000 1.4400 4.9600 1.5400 ;
      RECT 4.8700 0.7600 4.9600 1.4400 ;
      RECT 3.8850 0.6700 4.9600 0.7600 ;
      RECT 0.0450 0.4800 1.5200 0.5700 ;
      RECT 1.3050 0.4600 1.5200 0.4800 ;
      RECT 0.0450 1.8300 1.2300 1.9200 ;
      RECT 0.0450 1.3900 0.1700 1.8300 ;
      RECT 0.0450 0.7950 0.1350 1.3900 ;
      RECT 0.0450 0.5700 0.1700 0.7950 ;
  END
END CGENCON_X1P4M_A12TH

MACRO CGENCON_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 4.4750 1.9650 4.5850 2.0800 ;
        RECT 5.0100 1.9600 5.1200 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 1.2500 1.1700 1.3500 ;
        RECT 0.6200 1.0450 0.7550 1.2500 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END A

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6150 0.8750 4.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.1692 ;
  END CI

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9150 1.0500 1.6000 1.1500 ;
        RECT 1.5000 1.1500 1.6000 1.2500 ;
        RECT 1.5000 0.9500 1.6000 1.0500 ;
        RECT 1.5000 1.2500 1.8050 1.3500 ;
        RECT 1.5000 0.8400 1.7300 0.9500 ;
        RECT 1.7050 1.3500 1.8050 1.4600 ;
        RECT 1.7050 1.4600 2.2150 1.5600 ;
        RECT 2.1150 1.2300 2.2150 1.4600 ;
        RECT 2.1150 1.1200 2.4000 1.2300 ;
    END
    ANTENNAGATEAREA 0.2892 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.2900 0.3200 0.7100 0.3700 ;
        RECT 2.4050 0.3200 2.5050 0.6400 ;
        RECT 2.9150 0.3200 3.0250 0.5800 ;
    END
  END VSS

  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1200 1.6500 4.3100 1.7500 ;
        RECT 4.2100 1.7500 4.3100 1.7600 ;
        RECT 4.2100 1.7600 5.1500 1.8600 ;
        RECT 5.0500 0.5800 5.1500 1.7600 ;
        RECT 3.1200 0.4800 5.1500 0.5800 ;
        RECT 3.1200 0.4700 3.3350 0.4800 ;
    END
    ANTENNADIFFAREA 0.501375 ;
  END CON
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5200 0.5700 ;
      RECT 1.3050 0.4600 1.5200 0.4800 ;
      RECT 0.0450 1.8300 1.2300 1.9200 ;
      RECT 0.0450 1.3900 0.1700 1.8300 ;
      RECT 0.0450 0.7950 0.1350 1.3900 ;
      RECT 0.0450 0.5700 0.1700 0.7950 ;
      RECT 0.2600 0.6600 1.9900 0.7500 ;
      RECT 1.9000 0.7500 1.9900 1.1300 ;
      RECT 1.9000 1.1300 2.0100 1.3700 ;
      RECT 0.2600 1.6200 0.7300 1.7300 ;
      RECT 0.2600 1.1550 0.3500 1.6200 ;
      RECT 0.2300 0.9050 0.3500 1.1550 ;
      RECT 0.2600 0.7500 0.3500 0.9050 ;
      RECT 2.9750 1.9200 3.3950 1.9600 ;
      RECT 1.3250 1.8700 3.3950 1.9200 ;
      RECT 1.3250 1.8300 3.0650 1.8700 ;
      RECT 1.3250 1.7100 1.4150 1.8300 ;
      RECT 0.8300 1.6200 1.4150 1.7100 ;
      RECT 0.8300 1.5300 0.9400 1.6200 ;
      RECT 0.4400 1.4400 0.9400 1.5300 ;
      RECT 0.4400 0.8400 1.2800 0.9300 ;
      RECT 0.4400 0.9300 0.5300 1.4400 ;
      RECT 2.6700 1.2900 3.5950 1.3800 ;
      RECT 3.3400 1.2700 3.5950 1.2900 ;
      RECT 2.2900 0.7400 3.6050 0.7600 ;
      RECT 2.6600 0.6700 3.6050 0.7400 ;
      RECT 2.6700 1.3800 2.7600 1.5400 ;
      RECT 2.6700 0.8500 2.7600 1.2900 ;
      RECT 2.2900 0.7600 2.7600 0.8500 ;
      RECT 2.6600 0.4500 2.7700 0.6700 ;
      RECT 2.9100 1.4700 3.7850 1.5600 ;
      RECT 3.6950 1.2550 3.7850 1.4700 ;
      RECT 3.6950 1.1650 4.2750 1.2550 ;
      RECT 3.6950 0.9650 3.7850 1.1650 ;
      RECT 3.2350 0.8750 3.7850 0.9650 ;
      RECT 1.5250 1.6500 3.0000 1.7400 ;
      RECT 2.9100 1.5600 3.0000 1.6500 ;
      RECT 2.0900 0.6200 2.1800 0.9400 ;
      RECT 2.0900 0.5700 2.2850 0.6200 ;
      RECT 1.6100 0.4800 2.2850 0.5700 ;
      RECT 1.5250 1.5300 1.6150 1.6500 ;
      RECT 1.3000 1.4400 1.6150 1.5300 ;
      RECT 1.6100 0.4600 1.8200 0.4800 ;
      RECT 2.4900 1.0300 2.5800 1.6500 ;
      RECT 2.0900 0.9400 2.5800 1.0300 ;
      RECT 4.7250 1.5250 4.8850 1.6700 ;
      RECT 3.8850 1.4250 4.8850 1.5250 ;
      RECT 4.7250 1.3850 4.8850 1.4250 ;
      RECT 4.7250 1.2850 4.9600 1.3850 ;
      RECT 4.8700 0.7600 4.9600 1.2850 ;
      RECT 3.8850 0.6700 4.9600 0.7600 ;
  END
END CGENCON_X2M_A12TH

MACRO CGENI_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 1.3950 0.3200 1.4950 0.5800 ;
    END
  END VSS

  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7700 1.5500 1.4400 ;
        RECT 0.3200 1.4400 1.5500 1.5500 ;
        RECT 0.3050 0.6700 1.5500 0.7700 ;
        RECT 0.3200 1.5500 0.4900 1.7300 ;
    END
    ANTENNADIFFAREA 0.326 ;
  END CON

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8400 1.8900 1.0100 2.0800 ;
        RECT 1.3950 1.7800 1.4950 2.0800 ;
    END
  END VDD

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9450 0.3550 1.3500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5150 1.2500 1.3350 1.3500 ;
        RECT 0.5150 1.0100 0.6150 1.2500 ;
        RECT 1.2350 1.0050 1.3350 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7250 1.0450 1.1250 1.1500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.6300 1.6500 1.2700 1.7500 ;
      RECT 1.1000 1.7500 1.2700 1.9500 ;
      RECT 0.0950 1.8200 0.7300 1.9200 ;
      RECT 0.6300 1.7500 0.7300 1.8200 ;
      RECT 0.0950 1.5000 0.1950 1.8200 ;
      RECT 0.0950 0.4800 1.2850 0.5800 ;
      RECT 0.0950 0.5800 0.1950 0.8550 ;
  END
END CGENI_X1M_A12TH

MACRO CGENI_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.0450 1.8800 1.2150 2.0800 ;
        RECT 1.5650 1.8800 1.7350 2.0800 ;
        RECT 2.1200 1.7600 2.2200 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 1.0450 0.3200 1.2150 0.4950 ;
        RECT 1.5650 0.3200 1.7350 0.4950 ;
        RECT 2.1200 0.3200 2.2200 0.7150 ;
    END
  END VSS

  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4700 2.7550 1.5700 ;
        RECT 0.0800 1.5700 0.1800 1.8950 ;
        RECT 2.6200 1.5700 2.7550 1.8750 ;
        RECT 0.4800 1.4500 2.7550 1.4700 ;
        RECT 2.6650 0.8100 2.7550 1.4500 ;
        RECT 0.4800 0.7900 0.5800 1.4500 ;
        RECT 2.5850 0.4700 2.7550 0.8100 ;
        RECT 0.0450 0.6900 0.7600 0.7900 ;
        RECT 0.0450 0.4900 0.2150 0.6900 ;
    END
    ANTENNADIFFAREA 0.6318 ;
  END CON

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9350 1.0500 2.2800 1.1500 ;
        RECT 1.9350 0.9550 2.0350 1.0500 ;
        RECT 1.2200 0.8550 2.0350 0.9550 ;
        RECT 1.2200 0.9550 1.3200 1.0500 ;
        RECT 0.9300 1.0500 1.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2916 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.2500 2.5750 1.3500 ;
        RECT 1.4650 1.2000 1.8350 1.2500 ;
        RECT 2.4750 0.9400 2.5750 1.2500 ;
        RECT 0.6950 0.9150 0.7950 1.2500 ;
    END
    ANTENNAGATEAREA 0.2916 ;
  END A

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1850 1.2500 0.3900 1.3500 ;
        RECT 0.1850 0.9150 0.2850 1.2500 ;
    END
    ANTENNAGATEAREA 0.1458 ;
  END CI
  OBS
    LAYER M1 ;
      RECT 0.3050 1.6600 1.9950 1.7600 ;
      RECT 1.8250 1.7600 1.9950 1.9550 ;
      RECT 0.3050 1.7600 0.4750 1.9500 ;
      RECT 1.3050 1.7600 1.4750 1.9500 ;
      RECT 0.8500 0.6650 1.9950 0.7650 ;
      RECT 1.8250 0.4650 1.9950 0.6650 ;
      RECT 0.8500 0.5800 0.9500 0.6650 ;
      RECT 0.3050 0.4800 0.9500 0.5800 ;
      RECT 1.3050 0.4650 1.4750 0.6650 ;
  END
END CGENI_X1P4M_A12TH

MACRO CGENI_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.0450 1.8800 1.2150 2.0800 ;
        RECT 1.5650 1.8800 1.7350 2.0800 ;
        RECT 2.1200 1.7600 2.2200 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 2.1200 0.3200 2.2200 0.6100 ;
    END
  END VSS

  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.4500 2.7550 1.5500 ;
        RECT 0.0800 1.5500 0.1800 1.8950 ;
        RECT 2.6200 1.5500 2.7550 1.8750 ;
        RECT 2.6650 0.8100 2.7550 1.4500 ;
        RECT 0.4800 0.7900 0.5800 1.4500 ;
        RECT 2.5850 0.4700 2.7550 0.8100 ;
        RECT 0.0450 0.6900 0.7650 0.7900 ;
        RECT 0.0450 0.4900 0.2150 0.6900 ;
    END
    ANTENNADIFFAREA 0.8372 ;
  END CON

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9350 1.0500 2.2800 1.1500 ;
        RECT 1.9350 0.7900 2.0350 1.0500 ;
        RECT 1.2200 0.6900 2.0350 0.7900 ;
        RECT 1.2200 0.7900 1.3200 1.0500 ;
        RECT 1.0700 1.0500 1.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.3864 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.2500 2.5750 1.3500 ;
        RECT 1.4350 1.0750 1.5250 1.2500 ;
        RECT 2.4750 0.9400 2.5750 1.2500 ;
        RECT 0.6950 0.9150 0.7950 1.2500 ;
        RECT 1.4350 0.9750 1.7100 1.0750 ;
    END
    ANTENNAGATEAREA 0.3864 ;
  END A

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9100 0.3600 1.3600 ;
    END
    ANTENNAGATEAREA 0.1932 ;
  END CI
  OBS
    LAYER M1 ;
      RECT 0.3050 1.6450 1.9950 1.7450 ;
      RECT 1.8250 1.7450 1.9950 1.9550 ;
      RECT 0.3050 1.7450 0.4750 1.9500 ;
      RECT 1.3050 1.7450 1.4750 1.9500 ;
      RECT 0.3050 0.4800 2.0250 0.5800 ;
  END
END CGENI_X2M_A12TH

MACRO CGEN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.7950 1.8100 0.8950 2.0800 ;
        RECT 1.3300 1.7600 1.4300 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6550 0.8500 1.0600 0.9850 ;
    END
    ANTENNAGATEAREA 0.1812 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 1.2950 0.3200 1.4650 0.5150 ;
    END
  END VSS

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1750 0.8500 0.3500 1.2550 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END CI

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6450 0.8900 1.7500 1.3400 ;
        RECT 1.6100 1.3400 1.7500 1.4400 ;
        RECT 1.6100 0.7900 1.7500 0.8900 ;
        RECT 1.6100 1.4400 1.7100 1.8000 ;
        RECT 1.6100 0.4600 1.7100 0.7900 ;
    END
    ANTENNADIFFAREA 0.27625 ;
  END CO

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.2500 1.2550 1.3500 ;
        RECT 1.1650 0.8700 1.2550 1.2500 ;
        RECT 0.4450 0.8500 0.5550 1.2500 ;
    END
    ANTENNAGATEAREA 0.1812 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0750 1.6200 1.1900 1.7200 ;
      RECT 1.0200 1.7200 1.1900 1.9100 ;
      RECT 0.0750 1.7200 0.1750 1.9900 ;
      RECT 0.0700 0.5700 0.1900 0.7100 ;
      RECT 0.0700 0.4800 1.1900 0.5700 ;
      RECT 1.0100 0.4600 1.1900 0.4800 ;
      RECT 0.2800 1.4400 1.5200 1.5300 ;
      RECT 1.4300 0.7600 1.5200 1.4400 ;
      RECT 0.3000 0.6700 1.5200 0.7600 ;
  END
END CGEN_X1M_A12TH

MACRO CGEN_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.8950 1.8100 0.9950 2.0800 ;
        RECT 1.4300 1.7600 1.5300 2.0800 ;
        RECT 2.0000 1.7600 2.1000 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7400 0.8500 1.1900 0.9850 ;
    END
    ANTENNAGATEAREA 0.1812 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 1.3950 0.3200 1.5650 0.5150 ;
        RECT 1.9950 0.3200 2.0950 0.6050 ;
    END
  END VSS

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 0.8500 0.3500 1.2550 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END CI

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7100 1.4500 2.1450 1.5500 ;
        RECT 1.7100 1.5500 1.8100 1.9650 ;
        RECT 2.0550 0.9500 2.1450 1.4500 ;
        RECT 1.7100 0.8500 2.1450 0.9500 ;
        RECT 1.7100 0.5000 1.8100 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END CO

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.2500 1.3800 1.3500 ;
        RECT 1.2900 0.8700 1.3800 1.2500 ;
        RECT 0.4400 0.8500 0.5600 1.2500 ;
    END
    ANTENNAGATEAREA 0.1812 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0900 1.6200 1.2900 1.7200 ;
      RECT 1.1200 1.7200 1.2900 1.9100 ;
      RECT 0.0900 1.7200 0.1900 1.9900 ;
      RECT 0.0850 0.5700 0.2050 0.7100 ;
      RECT 0.0850 0.4800 1.2900 0.5700 ;
      RECT 1.1100 0.4600 1.2900 0.4800 ;
      RECT 1.4900 1.0500 1.8100 1.1500 ;
      RECT 0.2950 1.4400 1.5800 1.5300 ;
      RECT 1.4900 1.1500 1.5800 1.4400 ;
      RECT 1.4900 0.7600 1.5800 1.0500 ;
      RECT 0.3150 0.6700 1.5800 0.7600 ;
  END
END CGEN_X1P4M_A12TH

MACRO CGEN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.8950 1.8100 0.9950 2.0800 ;
        RECT 1.4300 1.7600 1.5300 2.0800 ;
        RECT 2.0000 1.7600 2.1000 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7350 0.8500 1.1900 0.9850 ;
    END
    ANTENNAGATEAREA 0.1812 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 1.3950 0.3200 1.5650 0.5150 ;
        RECT 1.9950 0.3200 2.0950 0.6050 ;
    END
  END VSS

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 0.8500 0.3500 1.2550 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END CI

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7100 1.2500 2.1450 1.3500 ;
        RECT 1.7100 1.3500 1.8100 1.7250 ;
        RECT 2.0550 0.9500 2.1450 1.2500 ;
        RECT 1.7100 0.8500 2.1450 0.9500 ;
        RECT 1.7100 0.4700 1.8100 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END CO

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.2500 1.3800 1.3500 ;
        RECT 1.2900 0.8700 1.3800 1.2500 ;
        RECT 0.4400 0.8500 0.5600 1.2500 ;
    END
    ANTENNAGATEAREA 0.1812 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0900 1.6200 1.2900 1.7200 ;
      RECT 1.1200 1.7200 1.2900 1.9100 ;
      RECT 0.0900 1.7200 0.1900 1.9900 ;
      RECT 0.0850 0.5700 0.2050 0.7100 ;
      RECT 0.0850 0.4800 1.2900 0.5700 ;
      RECT 1.1100 0.4600 1.2900 0.4800 ;
      RECT 1.4900 1.0500 1.8100 1.1500 ;
      RECT 0.2950 1.4400 1.5800 1.5300 ;
      RECT 1.4900 1.1500 1.5800 1.4400 ;
      RECT 1.4900 0.7600 1.5800 1.0500 ;
      RECT 0.3150 0.6700 1.5800 0.7600 ;
  END
END CGEN_X2M_A12TH

MACRO CMPR42_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 4.3850 2.0150 4.5550 2.0800 ;
        RECT 2.3700 1.8300 2.4700 2.0800 ;
        RECT 0.8600 1.8000 0.9600 2.0800 ;
        RECT 3.6450 1.7650 3.7450 2.0800 ;
        RECT 0.3350 1.7600 0.4350 2.0800 ;
        RECT 7.2050 1.7600 7.3050 2.0800 ;
        RECT 7.7250 1.7600 7.8250 2.0800 ;
        RECT 1.8500 1.6200 1.9500 2.0800 ;
    END
  END VDD

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1600 1.4500 4.4850 1.5500 ;
        RECT 4.1600 1.5500 4.2600 1.7200 ;
        RECT 4.1600 0.4450 4.2600 1.4500 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END SUM

  PIN ICI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8800 1.0500 7.6650 1.1500 ;
        RECT 5.8800 0.9850 5.9800 1.0500 ;
        RECT 7.5750 0.9200 7.6650 1.0500 ;
        RECT 4.8200 0.8950 5.9800 0.9850 ;
        RECT 4.8200 0.9850 4.9200 1.1050 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END ICI

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.3300 0.3200 0.4400 0.6400 ;
        RECT 0.8050 0.3200 1.0150 0.3650 ;
        RECT 1.8500 0.3200 1.9500 0.5800 ;
        RECT 6.2050 0.3200 6.3050 0.5800 ;
        RECT 7.1500 0.3200 7.3400 0.3750 ;
        RECT 7.7200 0.3200 7.8300 0.6300 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0800 0.8500 7.4250 0.9500 ;
        RECT 6.0800 0.8050 6.1800 0.8500 ;
        RECT 4.5900 0.7050 6.1800 0.8050 ;
        RECT 4.5900 0.8050 4.6900 1.1600 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END D

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0500 0.9000 8.1500 1.3000 ;
        RECT 7.9850 1.3000 8.1500 1.4000 ;
        RECT 7.9850 0.8000 8.1500 0.9000 ;
        RECT 7.9850 1.4000 8.0850 1.7600 ;
        RECT 7.9850 0.4350 8.0850 0.8000 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END CO

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5450 1.0500 2.1150 1.1500 ;
        RECT 2.0150 1.0000 2.1150 1.0500 ;
        RECT 2.0150 0.9000 3.1400 1.0000 ;
    END
    ANTENNAGATEAREA 0.201 ;
  END C

  PIN ICO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9100 0.1500 1.2900 ;
        RECT 0.0500 1.2900 0.1750 1.3900 ;
        RECT 0.0500 0.8100 0.1750 0.9100 ;
        RECT 0.0750 1.3900 0.1750 1.7750 ;
        RECT 0.0750 0.4500 0.1750 0.8100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END ICO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7200 1.0450 1.1250 1.1500 ;
        RECT 1.0150 0.9400 1.1250 1.0450 ;
        RECT 1.0150 0.8400 1.8500 0.9400 ;
        RECT 1.7500 0.8000 1.8500 0.8400 ;
        RECT 1.7500 0.7000 3.6100 0.8000 ;
        RECT 3.5100 0.8000 3.6100 1.1850 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.2500 2.3100 1.3500 ;
        RECT 2.2200 1.1900 2.3100 1.2500 ;
        RECT 1.2350 1.0300 1.3350 1.2500 ;
        RECT 0.4950 0.9850 0.5950 1.2500 ;
        RECT 2.2200 1.1000 3.3400 1.1900 ;
        RECT 3.2500 1.1900 3.3400 1.3700 ;
        RECT 3.2500 0.9150 3.3400 1.1000 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END A
  OBS
    LAYER M1 ;
      RECT 2.0750 1.6300 2.7650 1.7300 ;
      RECT 2.5950 1.7300 2.7650 1.9500 ;
      RECT 2.0750 1.7300 2.2450 1.9500 ;
      RECT 2.0500 0.4800 2.7650 0.5800 ;
      RECT 2.5600 0.4700 2.7650 0.4800 ;
      RECT 0.2650 1.4400 2.7650 1.5300 ;
      RECT 2.6750 1.3750 2.7650 1.4400 ;
      RECT 2.6750 1.2850 2.8900 1.3750 ;
      RECT 0.2650 0.8350 0.3550 1.4400 ;
      RECT 0.2650 0.7500 0.7500 0.8350 ;
      RECT 0.2650 0.7450 1.4950 0.7500 ;
      RECT 0.6600 0.6600 1.4950 0.7450 ;
      RECT 2.8900 1.5000 3.8000 1.5900 ;
      RECT 3.7100 1.1700 3.8000 1.5000 ;
      RECT 3.7100 0.9700 3.8500 1.1700 ;
      RECT 3.7100 0.5700 3.8000 0.9700 ;
      RECT 2.8550 0.4800 3.8000 0.5700 ;
      RECT 2.8900 1.5900 2.9900 1.9350 ;
      RECT 2.8550 0.4600 3.0400 0.4800 ;
      RECT 5.1600 1.3600 5.2500 1.7200 ;
      RECT 4.3500 1.2700 5.2500 1.3600 ;
      RECT 4.3500 0.4800 5.2900 0.5700 ;
      RECT 4.3500 0.5700 4.4400 1.2700 ;
      RECT 5.3800 1.5400 5.5500 1.7350 ;
      RECT 5.3800 1.4400 6.0800 1.5400 ;
      RECT 5.9100 1.5400 6.0800 1.7350 ;
      RECT 5.3800 0.4800 6.1050 0.5700 ;
      RECT 3.8900 1.8300 6.2150 1.9200 ;
      RECT 6.0150 1.9200 6.2150 1.9900 ;
      RECT 3.8900 1.4900 4.0300 1.8300 ;
      RECT 3.9400 0.8500 4.0300 1.4900 ;
      RECT 3.8900 0.4100 4.0300 0.8500 ;
      RECT 5.0150 1.9200 5.1850 1.9900 ;
      RECT 6.4650 1.5450 7.5650 1.6350 ;
      RECT 7.4650 1.6350 7.5650 1.9600 ;
      RECT 6.4650 1.6350 6.5650 1.9650 ;
      RECT 6.4700 0.5700 6.5600 0.7250 ;
      RECT 6.4700 0.4800 7.6250 0.5700 ;
      RECT 7.4050 0.4600 7.6250 0.4800 ;
      RECT 6.3000 1.3550 7.8550 1.4450 ;
      RECT 7.7650 1.1750 7.8550 1.3550 ;
      RECT 7.7650 1.0200 7.9350 1.1750 ;
      RECT 7.7650 0.8100 7.8550 1.0200 ;
      RECT 7.5300 0.7600 7.8550 0.8100 ;
      RECT 6.6700 0.7200 7.8550 0.7600 ;
      RECT 6.6700 0.6700 7.6200 0.7200 ;
      RECT 5.3650 1.1650 5.4550 1.2400 ;
      RECT 5.2200 1.0750 5.4550 1.1650 ;
      RECT 6.3000 1.3300 6.3900 1.3550 ;
      RECT 5.3650 1.2400 6.3900 1.3300 ;
      RECT 0.5650 1.6200 1.7350 1.7100 ;
      RECT 1.5650 1.7100 1.7350 1.9500 ;
      RECT 0.5650 1.7100 0.7350 1.9500 ;
      RECT 0.5400 0.4800 1.7550 0.5700 ;
  END
END CMPR42_X1M_A12TH

MACRO CMPR42_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6800 ;
        RECT 0.5900 0.3200 0.7000 0.6400 ;
        RECT 1.0600 0.3200 1.2700 0.3650 ;
        RECT 4.3050 0.3200 4.4050 0.5750 ;
        RECT 6.5900 0.3200 6.6900 0.5650 ;
        RECT 7.5300 0.3200 7.7200 0.3750 ;
        RECT 8.1000 0.3200 8.2100 0.6200 ;
        RECT 8.6250 0.3200 8.7250 0.6700 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.2500 2.7750 1.3500 ;
        RECT 2.6850 1.1900 2.7750 1.2500 ;
        RECT 1.4900 1.0500 1.5900 1.2500 ;
        RECT 0.7500 0.9850 0.8500 1.2500 ;
        RECT 2.6850 1.1000 3.5550 1.1900 ;
        RECT 3.4650 1.1900 3.5550 1.3700 ;
        RECT 3.4650 0.9150 3.5550 1.1000 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9750 1.0450 1.3900 1.1500 ;
        RECT 1.2800 0.9400 1.3900 1.0450 ;
        RECT 1.2800 0.8400 2.3650 0.9400 ;
        RECT 2.2650 0.8000 2.3650 0.8400 ;
        RECT 2.2650 0.7000 3.8000 0.8000 ;
        RECT 3.7000 0.8000 3.8000 1.1850 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END B

  PIN ICO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.4500 ;
        RECT 0.0500 1.4500 0.4350 1.5500 ;
        RECT 0.0500 0.8500 0.4350 0.9500 ;
        RECT 0.3350 1.5500 0.4350 1.9700 ;
        RECT 0.3350 0.4100 0.4350 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END ICO

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 4.2700 2.0150 4.4400 2.0800 ;
        RECT 4.7900 2.0150 4.9600 2.0800 ;
        RECT 2.0600 1.8600 2.1600 2.0800 ;
        RECT 2.5800 1.8300 2.6800 2.0800 ;
        RECT 1.1150 1.8000 1.2150 2.0800 ;
        RECT 3.8350 1.7650 3.9350 2.0800 ;
        RECT 0.0750 1.7600 0.1750 2.0800 ;
        RECT 0.5950 1.7600 0.6950 2.0800 ;
        RECT 7.5850 1.7600 7.6850 2.0800 ;
        RECT 8.1050 1.7600 8.2050 2.0800 ;
        RECT 8.6250 1.7600 8.7250 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8000 1.0500 2.5750 1.1500 ;
        RECT 2.4750 1.0000 2.5750 1.0500 ;
        RECT 2.4750 0.9000 3.3500 1.0000 ;
    END
    ANTENNAGATEAREA 0.201 ;
  END C

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9500 4.5500 1.2500 ;
        RECT 4.4500 1.2500 4.6650 1.3500 ;
        RECT 4.4500 0.8500 4.6650 0.9500 ;
        RECT 4.5650 1.3500 4.6650 1.7200 ;
        RECT 4.5650 0.5000 4.6650 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END SUM

  PIN ICI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2650 1.0500 8.0450 1.1500 ;
        RECT 6.2650 0.9850 6.3650 1.0500 ;
        RECT 7.9550 0.9200 8.0450 1.0500 ;
        RECT 5.1950 0.8950 6.3650 0.9850 ;
        RECT 5.1950 0.9850 5.2950 1.1050 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END ICI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4650 0.8500 7.8050 0.9500 ;
        RECT 6.4650 0.8050 6.5650 0.8500 ;
        RECT 4.9450 0.7050 6.5650 0.8050 ;
        RECT 4.9450 0.8050 5.0450 1.1600 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END D

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.6500 0.9500 8.7500 1.4500 ;
        RECT 8.3650 1.4500 8.7500 1.5500 ;
        RECT 8.3650 0.8500 8.7500 0.9500 ;
        RECT 8.3650 1.5500 8.4650 1.9700 ;
        RECT 8.3650 0.4100 8.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END CO
  OBS
    LAYER M1 ;
      RECT 1.8600 0.5700 1.9500 0.7300 ;
      RECT 0.7950 0.4800 1.9500 0.5700 ;
      RECT 0.8200 1.6200 2.0000 1.7100 ;
      RECT 0.8200 1.7100 0.9900 1.9500 ;
      RECT 2.2850 1.6300 2.9750 1.7300 ;
      RECT 2.8050 1.7300 2.9750 1.9500 ;
      RECT 2.2850 1.7300 2.4550 1.9500 ;
      RECT 2.2600 0.4800 2.9750 0.5800 ;
      RECT 2.7700 0.4700 2.9750 0.4800 ;
      RECT 0.5250 1.4400 2.9750 1.5300 ;
      RECT 2.8850 1.3750 2.9750 1.4400 ;
      RECT 2.8850 1.2850 3.0800 1.3750 ;
      RECT 0.5250 1.1450 0.6150 1.4400 ;
      RECT 0.2800 1.0550 0.6150 1.1450 ;
      RECT 0.5250 0.8350 0.6150 1.0550 ;
      RECT 0.5250 0.7500 1.0050 0.8350 ;
      RECT 0.5250 0.7450 1.7500 0.7500 ;
      RECT 0.9150 0.6600 1.7500 0.7450 ;
      RECT 3.1000 1.5000 3.9900 1.5900 ;
      RECT 3.9000 1.1700 3.9900 1.5000 ;
      RECT 3.9000 0.9700 4.0400 1.1700 ;
      RECT 3.9000 0.5700 3.9900 0.9700 ;
      RECT 3.0650 0.4800 3.9900 0.5700 ;
      RECT 3.1000 1.5900 3.2000 1.9300 ;
      RECT 3.0650 0.4600 3.2500 0.4800 ;
      RECT 5.5450 1.3600 5.6350 1.7200 ;
      RECT 4.7550 1.2700 5.6350 1.3600 ;
      RECT 4.7550 0.4800 5.6750 0.5700 ;
      RECT 4.7550 1.1550 4.8450 1.2700 ;
      RECT 4.6400 1.0450 4.8450 1.1550 ;
      RECT 4.7550 0.5700 4.8450 1.0450 ;
      RECT 5.7650 1.5400 5.9350 1.7350 ;
      RECT 5.7650 1.4400 6.4650 1.5400 ;
      RECT 6.2950 1.5400 6.4650 1.7350 ;
      RECT 5.7650 0.4800 6.4900 0.5700 ;
      RECT 4.0800 1.8300 6.6000 1.9200 ;
      RECT 6.4000 1.9200 6.6000 1.9900 ;
      RECT 4.0800 1.2900 4.2200 1.8300 ;
      RECT 4.1300 0.8500 4.2200 1.2900 ;
      RECT 4.0800 0.6750 4.2200 0.8500 ;
      RECT 5.4000 1.9200 5.5700 1.9900 ;
      RECT 6.8450 1.5450 7.9450 1.6350 ;
      RECT 7.8450 1.6350 7.9450 1.9650 ;
      RECT 6.8450 1.6350 6.9450 1.9900 ;
      RECT 6.8500 0.5700 6.9400 0.7250 ;
      RECT 6.8500 0.4800 8.0050 0.5700 ;
      RECT 7.7850 0.4600 8.0050 0.4800 ;
      RECT 8.1450 1.0500 8.4750 1.1500 ;
      RECT 7.0050 1.3550 8.2350 1.4450 ;
      RECT 8.1450 1.1500 8.2350 1.3550 ;
      RECT 8.1450 0.8100 8.2350 1.0500 ;
      RECT 7.9100 0.7600 8.2350 0.8100 ;
      RECT 7.0500 0.7200 8.2350 0.7600 ;
      RECT 7.0500 0.6700 8.0000 0.7200 ;
      RECT 5.7500 1.1650 5.8400 1.2400 ;
      RECT 5.6050 1.0750 5.8400 1.1650 ;
      RECT 7.0050 1.3300 7.0950 1.3550 ;
      RECT 5.7500 1.2400 7.0950 1.3300 ;
  END
END CMPR42_X1P4M_A12TH

MACRO CMPR42_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 4.2700 2.0150 4.4400 2.0800 ;
        RECT 4.7900 2.0150 4.9600 2.0800 ;
        RECT 2.0600 1.8600 2.1600 2.0800 ;
        RECT 2.5800 1.8300 2.6800 2.0800 ;
        RECT 1.1150 1.8000 1.2150 2.0800 ;
        RECT 3.8350 1.7650 3.9350 2.0800 ;
        RECT 0.0750 1.7600 0.1750 2.0800 ;
        RECT 0.5950 1.7600 0.6950 2.0800 ;
        RECT 7.5850 1.7600 7.6850 2.0800 ;
        RECT 8.1050 1.7600 8.2050 2.0800 ;
        RECT 8.6250 1.7600 8.7250 2.0800 ;
    END
  END VDD

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.6500 0.9500 8.7500 1.2500 ;
        RECT 8.3650 1.2500 8.7500 1.3500 ;
        RECT 8.3650 0.8500 8.7500 0.9500 ;
        RECT 8.3650 1.3500 8.4650 1.7700 ;
        RECT 8.3650 0.4350 8.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END CO

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4650 0.8500 7.8050 0.9500 ;
        RECT 6.4650 0.8050 6.5650 0.8500 ;
        RECT 4.9450 0.7050 6.5650 0.8050 ;
        RECT 4.9450 0.8050 5.0450 1.1600 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END D

  PIN ICI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2650 1.0500 8.0450 1.1500 ;
        RECT 6.2650 0.9850 6.3650 1.0500 ;
        RECT 7.9550 0.9200 8.0450 1.0500 ;
        RECT 5.1950 0.8950 6.3650 0.9850 ;
        RECT 5.1950 0.9850 5.2950 1.1050 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END ICI

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9500 4.5500 1.2500 ;
        RECT 4.4500 1.2500 4.6650 1.3500 ;
        RECT 4.4500 0.8500 4.6650 0.9500 ;
        RECT 4.5650 1.3500 4.6650 1.7200 ;
        RECT 4.5650 0.4450 4.6650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END SUM

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8000 1.0500 2.5750 1.1500 ;
        RECT 2.4750 1.0000 2.5750 1.0500 ;
        RECT 2.4750 0.9000 3.3500 1.0000 ;
    END
    ANTENNAGATEAREA 0.201 ;
  END C

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6400 ;
        RECT 0.5900 0.3200 0.7000 0.6400 ;
        RECT 1.0600 0.3200 1.2700 0.3650 ;
        RECT 4.3050 0.3200 4.4050 0.5750 ;
        RECT 6.5900 0.3200 6.6900 0.5650 ;
        RECT 7.5300 0.3200 7.7200 0.3750 ;
        RECT 8.1000 0.3200 8.2100 0.6200 ;
        RECT 8.6250 0.3200 8.7250 0.6200 ;
    END
  END VSS

  PIN ICO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.2500 ;
        RECT 0.0500 1.2500 0.4350 1.3500 ;
        RECT 0.0500 0.8500 0.4350 0.9500 ;
        RECT 0.3350 1.3500 0.4350 1.7750 ;
        RECT 0.3350 0.4500 0.4350 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END ICO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9750 1.0450 1.3900 1.1500 ;
        RECT 1.2800 0.9400 1.3900 1.0450 ;
        RECT 1.2800 0.8400 2.3650 0.9400 ;
        RECT 2.2650 0.8000 2.3650 0.8400 ;
        RECT 2.2650 0.7000 3.8000 0.8000 ;
        RECT 3.7000 0.8000 3.8000 1.1850 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.2500 2.7750 1.3500 ;
        RECT 2.6850 1.1900 2.7750 1.2500 ;
        RECT 1.4900 1.0500 1.5900 1.2500 ;
        RECT 0.7500 0.9850 0.8500 1.2500 ;
        RECT 2.6850 1.1000 3.5550 1.1900 ;
        RECT 3.4650 1.1900 3.5550 1.3700 ;
        RECT 3.4650 0.9150 3.5550 1.1000 ;
    END
    ANTENNAGATEAREA 0.2838 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.8600 0.5700 1.9500 0.7300 ;
      RECT 0.7950 0.4800 1.9500 0.5700 ;
      RECT 0.8200 1.6200 2.0000 1.7100 ;
      RECT 0.8200 1.7100 0.9900 1.9500 ;
      RECT 2.2850 1.6300 2.9750 1.7300 ;
      RECT 2.8050 1.7300 2.9750 1.9500 ;
      RECT 2.2850 1.7300 2.4550 1.9500 ;
      RECT 2.2600 0.4800 2.9750 0.5800 ;
      RECT 2.7700 0.4700 2.9750 0.4800 ;
      RECT 0.5250 1.4400 2.9750 1.5300 ;
      RECT 2.8850 1.3750 2.9750 1.4400 ;
      RECT 2.8850 1.2850 3.0800 1.3750 ;
      RECT 0.5250 1.1450 0.6150 1.4400 ;
      RECT 0.2800 1.0550 0.6150 1.1450 ;
      RECT 0.5250 0.8350 0.6150 1.0550 ;
      RECT 0.5250 0.7500 1.0050 0.8350 ;
      RECT 0.5250 0.7450 1.7500 0.7500 ;
      RECT 0.9150 0.6600 1.7500 0.7450 ;
      RECT 3.1000 1.5000 3.9900 1.5900 ;
      RECT 3.9000 1.1700 3.9900 1.5000 ;
      RECT 3.9000 0.9700 4.0400 1.1700 ;
      RECT 3.9000 0.5700 3.9900 0.9700 ;
      RECT 3.0650 0.4800 3.9900 0.5700 ;
      RECT 3.1000 1.5900 3.2000 1.9300 ;
      RECT 3.0650 0.4600 3.2500 0.4800 ;
      RECT 5.5450 1.3600 5.6350 1.7200 ;
      RECT 4.7550 1.2700 5.6350 1.3600 ;
      RECT 4.7550 0.4800 5.6750 0.5700 ;
      RECT 4.7550 1.1550 4.8450 1.2700 ;
      RECT 4.6400 1.0450 4.8450 1.1550 ;
      RECT 4.7550 0.5700 4.8450 1.0450 ;
      RECT 5.7650 1.5400 5.9350 1.7350 ;
      RECT 5.7650 1.4400 6.4650 1.5400 ;
      RECT 6.2950 1.5400 6.4650 1.7350 ;
      RECT 5.7650 0.4800 6.4900 0.5700 ;
      RECT 4.0800 1.8300 6.6000 1.9200 ;
      RECT 6.4000 1.9200 6.6000 1.9900 ;
      RECT 4.0800 1.2900 4.2200 1.8300 ;
      RECT 4.1300 0.8500 4.2200 1.2900 ;
      RECT 4.0800 0.6750 4.2200 0.8500 ;
      RECT 5.4000 1.9200 5.5700 1.9900 ;
      RECT 6.8450 1.5450 7.9450 1.6350 ;
      RECT 7.8450 1.6350 7.9450 1.9650 ;
      RECT 6.8450 1.6350 6.9450 1.9900 ;
      RECT 6.8500 0.5700 6.9400 0.7250 ;
      RECT 6.8500 0.4800 8.0050 0.5700 ;
      RECT 7.7850 0.4600 8.0050 0.4800 ;
      RECT 8.1450 1.0500 8.4750 1.1500 ;
      RECT 7.0050 1.3550 8.2350 1.4450 ;
      RECT 8.1450 1.1500 8.2350 1.3550 ;
      RECT 8.1450 0.8100 8.2350 1.0500 ;
      RECT 7.9100 0.7600 8.2350 0.8100 ;
      RECT 7.0500 0.7200 8.2350 0.7600 ;
      RECT 7.0500 0.6700 8.0000 0.7200 ;
      RECT 5.7500 1.1650 5.8400 1.2400 ;
      RECT 5.6050 1.0750 5.8400 1.1650 ;
      RECT 7.0050 1.3300 7.0950 1.3550 ;
      RECT 5.7500 1.2400 7.0950 1.3300 ;
  END
END CMPR42_X2M_A12TH

MACRO DFFNQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 3.0050 0.3200 3.0950 0.7050 ;
        RECT 3.7300 0.3200 3.9000 0.5250 ;
    END
  END VSS

  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6400 1.0500 3.7500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END CKN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7350 0.5500 1.1900 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.9350 4.1500 1.3400 ;
        RECT 3.9850 1.3400 4.1500 1.7750 ;
        RECT 4.0300 0.5050 4.1500 0.9350 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7050 0.6850 0.7950 1.6950 ;
      RECT 1.0850 1.5250 1.4750 1.6150 ;
      RECT 1.3850 0.9300 1.4750 1.5250 ;
      RECT 1.3850 0.8400 1.7900 0.9300 ;
      RECT 1.7000 0.9300 1.7900 1.0500 ;
      RECT 1.3850 0.7500 1.4750 0.8400 ;
      RECT 1.0850 0.6600 1.4750 0.7500 ;
      RECT 1.9500 1.5400 2.1200 1.7400 ;
      RECT 1.9000 1.4500 2.1200 1.5400 ;
      RECT 1.9000 1.2300 1.9900 1.4500 ;
      RECT 1.5650 1.1400 1.9900 1.2300 ;
      RECT 1.9000 0.7500 1.9900 1.1400 ;
      RECT 1.9000 0.6600 2.1200 0.7500 ;
      RECT 2.2350 0.7750 2.6950 0.8650 ;
      RECT 2.2350 0.5700 2.3250 0.7750 ;
      RECT 0.0750 0.4800 2.3250 0.5700 ;
      RECT 0.8850 0.5700 0.9750 1.1950 ;
      RECT 0.0750 0.5700 0.1700 1.6850 ;
      RECT 2.7850 0.7950 3.1450 0.8850 ;
      RECT 3.0550 0.8850 3.1450 1.0050 ;
      RECT 2.3900 1.3250 2.4800 1.7200 ;
      RECT 2.3900 1.2350 2.8750 1.3250 ;
      RECT 2.7850 0.8850 2.8750 1.2350 ;
      RECT 2.7850 0.6400 2.8750 0.7950 ;
      RECT 2.4150 0.5500 2.8750 0.6400 ;
      RECT 0.2850 1.8300 3.5300 1.9200 ;
      RECT 3.4400 1.8000 3.5300 1.8300 ;
      RECT 0.8850 1.4150 0.9750 1.8300 ;
      RECT 2.2100 1.1700 2.3000 1.8300 ;
      RECT 3.4400 1.7000 3.6350 1.8000 ;
      RECT 0.8850 1.3250 1.2750 1.4150 ;
      RECT 2.1000 1.1250 2.3000 1.1700 ;
      RECT 3.4400 0.9050 3.5300 1.7000 ;
      RECT 1.1850 0.8650 1.2750 1.3250 ;
      RECT 2.1000 1.0350 2.6900 1.1250 ;
      RECT 3.4400 0.8150 3.6150 0.9050 ;
      RECT 2.1000 0.9600 2.1900 1.0350 ;
      RECT 0.2850 1.2600 0.3750 1.8300 ;
      RECT 3.2350 0.6250 3.9400 0.7150 ;
      RECT 3.8500 0.7150 3.9400 1.2150 ;
      RECT 3.2350 1.5050 3.3250 1.6350 ;
      RECT 2.7450 1.4150 3.3250 1.5050 ;
      RECT 3.2350 0.7150 3.3250 1.4150 ;
      RECT 3.2350 0.5050 3.3550 0.6250 ;
  END
END DFFNQ_X1M_A12TH

MACRO BUF_X0P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.7050 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8000 0.3600 1.1900 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7200 0.7500 1.3600 ;
        RECT 0.6300 1.3600 0.7500 1.8000 ;
        RECT 0.6250 0.5100 0.7500 0.7200 ;
    END
    ANTENNADIFFAREA 0.1552 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3650 1.5850 0.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.3000 0.5400 1.3900 ;
      RECT 0.4500 1.1000 0.5400 1.3000 ;
      RECT 0.0500 1.3900 0.1750 1.5500 ;
      RECT 0.0500 0.7200 0.1400 1.3000 ;
      RECT 0.0500 0.5300 0.1700 0.7200 ;
  END
END BUF_X0P7B_A12TH

MACRO BUF_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.7000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.5550 1.2200 ;
    END
    ANTENNAGATEAREA 0.0222 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7000 0.1500 1.5600 ;
        RECT 0.0500 1.5600 0.1700 1.9700 ;
        RECT 0.0500 0.5100 0.1750 0.7000 ;
    END
    ANTENNADIFFAREA 0.1848 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3350 1.7600 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6300 1.4700 0.7550 1.7150 ;
      RECT 0.2400 1.3800 0.7550 1.4700 ;
      RECT 0.6650 0.7200 0.7550 1.3800 ;
      RECT 0.6250 0.5300 0.7550 0.7200 ;
      RECT 0.2400 1.2050 0.3300 1.3800 ;
  END
END BUF_X0P7M_A12TH

MACRO BUF_X0P8B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3300 0.3200 0.5000 0.7000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8100 0.3600 1.1950 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.7000 0.7500 1.4800 ;
        RECT 0.6300 1.4800 0.7500 1.9100 ;
        RECT 0.6300 0.4900 0.7500 0.7000 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3650 1.7400 0.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0700 1.3050 0.5600 1.3950 ;
      RECT 0.4700 1.1050 0.5600 1.3050 ;
      RECT 0.0700 1.3950 0.1800 1.6300 ;
      RECT 0.0700 0.7400 0.1600 1.3050 ;
      RECT 0.0700 0.5500 0.1700 0.7400 ;
  END
END BUF_X0P8B_A12TH

MACRO BUF_X0P8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.7900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9000 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8100 0.1500 1.6600 ;
        RECT 0.0500 1.6600 0.1750 1.8700 ;
        RECT 0.0500 0.4300 0.1700 0.8100 ;
    END
    ANTENNADIFFAREA 0.2184 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3350 1.7600 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6250 1.5700 0.7500 1.6700 ;
      RECT 0.2400 1.4800 0.7500 1.5700 ;
      RECT 0.6600 0.7900 0.7500 1.4800 ;
      RECT 0.6250 0.6000 0.7500 0.7900 ;
      RECT 0.2400 1.1650 0.3300 1.4800 ;
  END
END BUF_X0P8M_A12TH

MACRO BUF_X11B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.7300 ;
        RECT 0.8650 0.3200 1.0350 0.7300 ;
        RECT 1.3850 0.3200 1.5550 0.7300 ;
        RECT 1.9050 0.3200 2.0750 0.7300 ;
        RECT 2.4250 0.3200 2.5950 0.7300 ;
        RECT 2.9450 0.3200 3.1150 0.7300 ;
        RECT 3.4650 0.3200 3.6350 0.7300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.3850 1.7700 0.4750 2.0800 ;
        RECT 0.9050 1.7700 0.9950 2.0800 ;
        RECT 1.4250 1.7700 1.5150 2.0800 ;
        RECT 1.9450 1.7700 2.0350 2.0800 ;
        RECT 2.4650 1.7700 2.5550 2.0800 ;
        RECT 2.9850 1.7700 3.0750 2.0800 ;
        RECT 3.5050 1.7700 3.5950 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7850 1.1500 ;
    END
    ANTENNAGATEAREA 0.2457 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1650 1.4200 3.8550 1.5800 ;
        RECT 1.1650 1.5800 1.2550 1.8500 ;
        RECT 1.6850 1.5800 1.7750 1.8500 ;
        RECT 2.2050 1.5800 2.2950 1.8500 ;
        RECT 2.7250 1.5800 2.8150 1.8500 ;
        RECT 3.2450 1.5800 3.3350 1.8500 ;
        RECT 3.7650 1.5800 3.8550 1.8500 ;
        RECT 3.4200 0.9800 3.5800 1.4200 ;
        RECT 1.1650 0.8200 3.8550 0.9800 ;
        RECT 1.1650 0.4500 1.2550 0.8200 ;
        RECT 1.6850 0.4500 1.7750 0.8200 ;
        RECT 2.2050 0.4500 2.2950 0.8200 ;
        RECT 2.7250 0.4500 2.8150 0.8200 ;
        RECT 3.2450 0.4500 3.3350 0.8200 ;
        RECT 3.7650 0.4500 3.8550 0.8200 ;
    END
    ANTENNADIFFAREA 1.644825 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.9200 1.0700 3.0750 1.1600 ;
      RECT 0.1250 1.3700 0.2150 1.7200 ;
      RECT 0.1250 0.4600 0.2150 0.8300 ;
      RECT 0.6450 1.3700 0.7350 1.7200 ;
      RECT 0.6450 0.4550 0.7350 0.8300 ;
      RECT 0.1250 1.2800 1.0100 1.3700 ;
      RECT 0.9200 1.1600 1.0100 1.2800 ;
      RECT 0.9200 0.9200 1.0100 1.0700 ;
      RECT 0.1250 0.8300 1.0100 0.9200 ;
  END
END BUF_X11B_A12TH

MACRO BUF_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3850 0.3200 0.4750 0.6300 ;
        RECT 0.9050 0.3200 0.9950 0.6300 ;
        RECT 1.4250 0.3200 1.5150 0.6300 ;
        RECT 1.9450 0.3200 2.0350 0.6300 ;
        RECT 2.4650 0.3200 2.5550 0.6300 ;
        RECT 2.9850 0.3200 3.0750 0.6300 ;
        RECT 3.5050 0.3200 3.5950 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.3850 1.7700 0.4750 2.0800 ;
        RECT 0.9050 1.7700 0.9950 2.0800 ;
        RECT 1.4250 1.7700 1.5150 2.0800 ;
        RECT 1.9450 1.7700 2.0350 2.0800 ;
        RECT 2.4650 1.7700 2.5550 2.0800 ;
        RECT 2.9850 1.7700 3.0750 2.0800 ;
        RECT 3.5050 1.7700 3.5950 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1650 1.4200 3.8550 1.5800 ;
        RECT 1.1650 1.5800 1.2550 1.8500 ;
        RECT 1.6850 1.5800 1.7750 1.8500 ;
        RECT 2.2050 1.5800 2.2950 1.8500 ;
        RECT 2.7250 1.5800 2.8150 1.8500 ;
        RECT 3.2450 1.5800 3.3350 1.8500 ;
        RECT 3.7650 1.5800 3.8550 1.8500 ;
        RECT 3.4200 0.9800 3.5800 1.4200 ;
        RECT 1.1650 0.8200 3.8550 0.9800 ;
        RECT 1.1650 0.4850 1.2550 0.8200 ;
        RECT 1.6850 0.4850 1.7750 0.8200 ;
        RECT 2.2050 0.4850 2.2950 0.8200 ;
        RECT 2.7250 0.4850 2.8150 0.8200 ;
        RECT 3.2450 0.4850 3.3350 0.8200 ;
        RECT 3.7650 0.4850 3.8550 0.8200 ;
    END
    ANTENNADIFFAREA 1.958125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2750 1.0500 0.7850 1.1500 ;
    END
    ANTENNAGATEAREA 0.2925 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.9200 1.0700 3.1300 1.1600 ;
      RECT 0.6450 1.3700 0.7350 1.7200 ;
      RECT 0.6450 0.4850 0.7350 0.8300 ;
      RECT 0.1250 1.2800 1.0100 1.3700 ;
      RECT 0.9200 1.1600 1.0100 1.2800 ;
      RECT 0.9200 0.9200 1.0100 1.0700 ;
      RECT 0.1250 0.8300 1.0100 0.9200 ;
      RECT 0.1250 1.3700 0.2150 1.7200 ;
      RECT 0.1250 0.4850 0.2150 0.8300 ;
  END
END BUF_X11M_A12TH

MACRO BUF_X13B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.1300 0.3200 0.2200 0.9150 ;
        RECT 0.6500 0.3200 0.7400 0.7150 ;
        RECT 1.1700 0.3200 1.2600 0.7150 ;
        RECT 1.7050 0.3200 1.7950 0.6700 ;
        RECT 2.2250 0.3200 2.3150 0.6700 ;
        RECT 2.7450 0.3200 2.8350 0.6700 ;
        RECT 3.2650 0.3200 3.3550 0.6700 ;
        RECT 3.7850 0.3200 3.8750 0.6700 ;
        RECT 4.3050 0.3200 4.3950 0.6700 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2950 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2952 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.4100 4.6550 1.5900 ;
        RECT 1.4450 1.5900 1.5350 1.8800 ;
        RECT 1.9650 1.5900 2.0550 1.8800 ;
        RECT 2.4850 1.5900 2.5750 1.8800 ;
        RECT 3.0050 1.5900 3.0950 1.8800 ;
        RECT 3.5250 1.5900 3.6150 1.8800 ;
        RECT 4.0450 1.5900 4.1350 1.8800 ;
        RECT 4.5650 1.5900 4.6550 1.8800 ;
        RECT 4.0200 0.9900 4.1800 1.4100 ;
        RECT 1.4450 0.8100 4.6550 0.9900 ;
        RECT 1.4450 0.4950 1.5350 0.8100 ;
        RECT 1.9650 0.4950 2.0550 0.8100 ;
        RECT 2.4850 0.4950 2.5750 0.8100 ;
        RECT 3.0050 0.4950 3.0950 0.8100 ;
        RECT 3.5250 0.4950 3.6150 0.8100 ;
        RECT 4.0450 0.4950 4.1350 0.8100 ;
        RECT 4.5650 0.4950 4.6550 0.8100 ;
    END
    ANTENNADIFFAREA 1.917825 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 1.7050 1.7700 1.7950 2.0800 ;
        RECT 2.2250 1.7700 2.3150 2.0800 ;
        RECT 2.7450 1.7700 2.8350 2.0800 ;
        RECT 3.2650 1.7700 3.3550 2.0800 ;
        RECT 3.7850 1.7700 3.8750 2.0800 ;
        RECT 4.3050 1.7700 4.3950 2.0800 ;
        RECT 0.1300 1.6800 0.2200 2.0800 ;
        RECT 0.6500 1.6800 0.7400 2.0800 ;
        RECT 1.1850 1.6800 1.2750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.2000 1.0800 3.6950 1.1700 ;
      RECT 0.3900 1.3700 0.4800 1.7200 ;
      RECT 0.3900 0.4850 0.4800 0.8300 ;
      RECT 0.9100 1.3700 1.0000 1.7200 ;
      RECT 0.9100 0.4850 1.0000 0.8300 ;
      RECT 0.3900 1.2800 1.2900 1.3700 ;
      RECT 1.2000 1.1700 1.2900 1.2800 ;
      RECT 1.2000 0.9200 1.2900 1.0800 ;
      RECT 0.3900 0.8300 1.2900 0.9200 ;
  END
END BUF_X13B_A12TH

MACRO BUF_X13M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.1300 0.3200 0.2200 0.7100 ;
        RECT 0.6500 0.3200 0.7400 0.7100 ;
        RECT 1.1800 0.3200 1.2700 0.7100 ;
        RECT 1.7050 0.3200 1.7950 0.6300 ;
        RECT 2.2250 0.3200 2.3150 0.6300 ;
        RECT 2.7450 0.3200 2.8350 0.6300 ;
        RECT 3.2650 0.3200 3.3550 0.6300 ;
        RECT 3.7850 0.3200 3.8750 0.6300 ;
        RECT 4.3050 0.3200 4.3950 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 1.7050 1.7700 1.7950 2.0800 ;
        RECT 2.2250 1.7700 2.3150 2.0800 ;
        RECT 2.7450 1.7700 2.8350 2.0800 ;
        RECT 3.2650 1.7700 3.3550 2.0800 ;
        RECT 3.7850 1.7700 3.8750 2.0800 ;
        RECT 4.3050 1.7700 4.3950 2.0800 ;
        RECT 0.1300 1.6650 0.2200 2.0800 ;
        RECT 0.6500 1.6650 0.7400 2.0800 ;
        RECT 1.1850 1.6650 1.2750 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.4100 4.6550 1.5900 ;
        RECT 1.4450 1.5900 1.5350 1.8400 ;
        RECT 1.9650 1.5900 2.0550 1.8400 ;
        RECT 2.4850 1.5900 2.5750 1.8400 ;
        RECT 3.0050 1.5900 3.0950 1.8400 ;
        RECT 3.5250 1.5900 3.6150 1.8400 ;
        RECT 4.0450 1.5900 4.1350 1.8400 ;
        RECT 4.5650 1.5900 4.6550 1.8400 ;
        RECT 4.4200 0.9900 4.5800 1.4100 ;
        RECT 1.4450 0.8100 4.6550 0.9900 ;
        RECT 1.4450 0.4850 1.5350 0.8100 ;
        RECT 1.9650 0.4850 2.0550 0.8100 ;
        RECT 2.4850 0.4850 2.5750 0.8100 ;
        RECT 3.0050 0.4850 3.0950 0.8100 ;
        RECT 3.5250 0.4850 3.6150 0.8100 ;
        RECT 4.0450 0.4850 4.1350 0.8100 ;
        RECT 4.5650 0.4850 4.6550 0.8100 ;
    END
    ANTENNADIFFAREA 2.283125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.0500 0.9950 1.1500 ;
    END
    ANTENNAGATEAREA 0.3456 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.2350 1.0800 3.6800 1.1700 ;
      RECT 0.3900 1.3700 0.4800 1.7200 ;
      RECT 0.3900 0.5000 0.4800 0.8300 ;
      RECT 0.9100 1.3700 1.0000 1.7200 ;
      RECT 0.9100 0.5000 1.0000 0.8300 ;
      RECT 0.3900 1.2800 1.3250 1.3700 ;
      RECT 1.2350 1.1700 1.3250 1.2800 ;
      RECT 1.2350 0.9200 1.3250 1.0800 ;
      RECT 0.3900 0.8300 1.3250 0.9200 ;
  END
END BUF_X13M_A12TH

MACRO BUF_X16B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3950 0.3200 0.4850 0.6950 ;
        RECT 0.9150 0.3200 1.0050 0.6950 ;
        RECT 1.4500 0.3200 1.5400 0.6950 ;
        RECT 1.9300 0.3200 2.1000 0.6750 ;
        RECT 2.4500 0.3200 2.6200 0.6750 ;
        RECT 2.9700 0.3200 3.1400 0.6750 ;
        RECT 3.4900 0.3200 3.6600 0.6750 ;
        RECT 4.0100 0.3200 4.1800 0.6750 ;
        RECT 4.5300 0.3200 4.7000 0.6750 ;
        RECT 5.0500 0.3200 5.2200 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 1.9700 1.7700 2.0600 2.0800 ;
        RECT 2.4900 1.7700 2.5800 2.0800 ;
        RECT 3.0100 1.7700 3.1000 2.0800 ;
        RECT 3.5300 1.7700 3.6200 2.0800 ;
        RECT 4.0500 1.7700 4.1400 2.0800 ;
        RECT 4.5700 1.7700 4.6600 2.0800 ;
        RECT 5.0900 1.7700 5.1800 2.0800 ;
        RECT 5.6100 1.7700 5.7000 2.0800 ;
        RECT 0.3950 1.6750 0.4850 2.0800 ;
        RECT 0.9150 1.6750 1.0050 2.0800 ;
        RECT 1.4350 1.6750 1.5250 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7100 1.3900 5.4400 1.6100 ;
        RECT 1.7100 1.6100 1.8000 1.8200 ;
        RECT 2.2300 1.6100 2.3200 1.8200 ;
        RECT 2.7500 1.6100 2.8400 1.8200 ;
        RECT 3.2700 1.6100 3.3600 1.8200 ;
        RECT 3.7900 1.6100 3.8800 1.8200 ;
        RECT 4.3100 1.6100 4.4000 1.8200 ;
        RECT 4.8300 1.6100 4.9200 1.8200 ;
        RECT 5.3500 1.6100 5.4400 1.8200 ;
        RECT 4.9900 0.9900 5.2100 1.3900 ;
        RECT 1.7100 0.7700 5.2100 0.9900 ;
        RECT 4.8300 0.5000 4.9200 0.7700 ;
        RECT 1.7100 0.4800 1.8000 0.7700 ;
        RECT 2.2250 0.4800 2.3250 0.7700 ;
        RECT 2.7450 0.4800 2.8450 0.7700 ;
        RECT 3.2650 0.4800 3.3650 0.7700 ;
        RECT 3.7850 0.4800 3.8850 0.7700 ;
        RECT 4.3050 0.4800 4.4050 0.7700 ;
    END
    ANTENNADIFFAREA 2.184 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4200 1.0500 1.2300 1.1500 ;
    END
    ANTENNAGATEAREA 0.366 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.4650 1.1000 4.5250 1.1900 ;
      RECT 0.1350 1.3700 0.2250 1.7200 ;
      RECT 0.1350 0.4600 0.2250 0.8300 ;
      RECT 0.6550 1.3700 0.7450 1.7200 ;
      RECT 0.6550 0.4600 0.7450 0.8300 ;
      RECT 1.1750 1.3700 1.2650 1.7200 ;
      RECT 1.1750 0.4600 1.2650 0.8300 ;
      RECT 0.1350 1.2800 1.5550 1.3700 ;
      RECT 1.4650 1.1900 1.5550 1.2800 ;
      RECT 1.4650 0.9200 1.5550 1.1000 ;
      RECT 0.1350 0.8300 1.5550 0.9200 ;
  END
END BUF_X16B_A12TH

MACRO BUF_X16M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3950 0.3200 0.4850 0.7100 ;
        RECT 0.9150 0.3200 1.0050 0.7100 ;
        RECT 1.4350 0.3200 1.5250 0.7100 ;
        RECT 1.9700 0.3200 2.0600 0.6300 ;
        RECT 2.4900 0.3200 2.5800 0.6300 ;
        RECT 3.0100 0.3200 3.1000 0.6300 ;
        RECT 3.5300 0.3200 3.6200 0.6300 ;
        RECT 4.0500 0.3200 4.1400 0.6300 ;
        RECT 4.5700 0.3200 4.6600 0.6300 ;
        RECT 5.0900 0.3200 5.1800 0.6300 ;
        RECT 5.6100 0.3200 5.7000 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 1.9700 1.7700 2.0600 2.0800 ;
        RECT 2.4900 1.7700 2.5800 2.0800 ;
        RECT 3.0100 1.7700 3.1000 2.0800 ;
        RECT 3.5300 1.7700 3.6200 2.0800 ;
        RECT 4.0500 1.7700 4.1400 2.0800 ;
        RECT 4.5700 1.7700 4.6600 2.0800 ;
        RECT 5.0900 1.7700 5.1800 2.0800 ;
        RECT 5.6100 1.7700 5.7000 2.0800 ;
        RECT 0.3950 1.6600 0.4850 2.0800 ;
        RECT 0.9150 1.6600 1.0050 2.0800 ;
        RECT 1.4350 1.6600 1.5250 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4200 1.0500 1.2300 1.1500 ;
    END
    ANTENNAGATEAREA 0.429 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7100 1.3900 5.4400 1.6100 ;
        RECT 1.7100 1.6100 1.8000 1.8200 ;
        RECT 2.2300 1.6100 2.3200 1.8200 ;
        RECT 2.7500 1.6100 2.8400 1.8200 ;
        RECT 3.2700 1.6100 3.3600 1.8200 ;
        RECT 3.7900 1.6100 3.8800 1.8200 ;
        RECT 4.3100 1.6100 4.4000 1.8200 ;
        RECT 4.8300 1.6100 4.9200 1.8200 ;
        RECT 5.3500 1.6100 5.4400 1.8200 ;
        RECT 5.1900 0.9900 5.4400 1.3900 ;
        RECT 1.7100 0.7700 5.4400 0.9900 ;
        RECT 1.7100 0.4850 1.8000 0.7700 ;
        RECT 2.2300 0.4850 2.3200 0.7700 ;
        RECT 2.7500 0.4850 2.8400 0.7700 ;
        RECT 3.2700 0.4850 3.3600 0.7700 ;
        RECT 3.7900 0.4850 3.8800 0.7700 ;
        RECT 4.3100 0.4850 4.4000 0.7700 ;
        RECT 4.8300 0.4850 4.9200 0.7700 ;
        RECT 5.3500 0.4850 5.4400 0.7700 ;
    END
    ANTENNADIFFAREA 2.6 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.4650 1.1000 4.7900 1.1900 ;
      RECT 0.1350 1.3700 0.2250 1.7200 ;
      RECT 0.1350 0.4850 0.2250 0.8300 ;
      RECT 0.6550 1.3700 0.7450 1.7200 ;
      RECT 0.6550 0.4850 0.7450 0.8300 ;
      RECT 1.1750 1.3700 1.2650 1.7200 ;
      RECT 1.1750 0.4850 1.2650 0.8300 ;
      RECT 0.1350 1.2800 1.5550 1.3700 ;
      RECT 1.4650 1.1900 1.5550 1.2800 ;
      RECT 1.4650 0.9200 1.5550 1.1000 ;
      RECT 0.1350 0.8300 1.5550 0.9200 ;
  END
END BUF_X16M_A12TH

MACRO BUF_X1B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3000 0.3200 0.4700 0.6700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6750 0.1500 1.5250 ;
        RECT 0.0500 1.5250 0.1750 1.9350 ;
        RECT 0.0500 0.4650 0.1700 0.6750 ;
    END
    ANTENNADIFFAREA 0.2184 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.5600 1.2000 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3350 1.7700 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6250 1.4350 0.7400 1.5550 ;
      RECT 0.2400 1.3450 0.7400 1.4350 ;
      RECT 0.6500 0.7250 0.7400 1.3450 ;
      RECT 0.6300 0.4950 0.7400 0.7250 ;
      RECT 0.2400 0.9800 0.3300 1.3450 ;
  END
END BUF_X1B_A12TH

MACRO BUF_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9100 0.7500 1.5850 ;
        RECT 0.6300 1.5850 0.7500 1.9550 ;
        RECT 0.6300 0.5000 0.7500 0.9100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 1.0000 0.3500 1.1000 ;
        RECT 0.2500 1.1000 0.3500 1.3050 ;
    END
    ANTENNAGATEAREA 0.0294 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3650 1.7800 0.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5000 0.5400 1.5900 ;
      RECT 0.4500 0.9000 0.5400 1.5000 ;
      RECT 0.0800 0.8100 0.5400 0.9000 ;
      RECT 0.0800 1.4050 0.1700 1.5000 ;
      RECT 0.0800 0.7050 0.1700 0.8100 ;
  END
END BUF_X1M_A12TH

MACRO BUF_X1P2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4500 0.3200 0.6200 0.6700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.7300 1.2500 1.1500 1.3500 ;
        RECT 0.7450 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.3500 0.8200 1.7150 ;
        RECT 0.7450 0.4600 0.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.2079 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9650 0.3500 1.3500 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4300 1.6700 0.6000 2.0800 ;
        RECT 0.9900 1.4400 1.0800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0600 0.9150 1.1500 ;
      RECT 0.0750 1.4800 0.5500 1.5700 ;
      RECT 0.4600 1.1500 0.5500 1.4800 ;
      RECT 0.4600 0.8500 0.5500 1.0600 ;
      RECT 0.0750 0.7600 0.5500 0.8500 ;
  END
END BUF_X1P2B_A12TH

MACRO BUF_X1P2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.7050 ;
        RECT 0.9900 0.3200 1.0800 0.7050 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4700 1.6900 0.5600 2.0800 ;
        RECT 0.9900 1.4700 1.0800 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0348 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.7300 1.2500 1.1500 1.3500 ;
        RECT 0.7250 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.3500 0.8200 1.7900 ;
        RECT 0.7250 0.4850 0.8250 0.8500 ;
    END
    ANTENNADIFFAREA 0.193 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.5300 1.0600 0.9400 1.1500 ;
      RECT 0.0750 1.4800 0.6200 1.5700 ;
      RECT 0.5300 1.1500 0.6200 1.4800 ;
      RECT 0.5300 0.9150 0.6200 1.0600 ;
      RECT 0.1350 0.8250 0.6200 0.9150 ;
      RECT 0.1350 0.7050 0.2250 0.8250 ;
  END
END BUF_X1P2M_A12TH

MACRO BUF_X1P4B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4900 0.3200 0.5800 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.4500 ;
        RECT 0.7300 1.4500 1.1500 1.5500 ;
        RECT 0.7450 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.5500 0.8200 1.8800 ;
        RECT 0.7450 0.5200 0.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.26225 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.0100 0.3550 1.3700 ;
    END
    ANTENNAGATEAREA 0.0351 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.9900 1.6650 1.0800 2.0800 ;
        RECT 0.4700 1.6600 0.5600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4650 1.1750 0.9300 1.2650 ;
      RECT 0.0950 1.4800 0.5550 1.5700 ;
      RECT 0.4650 1.2650 0.5550 1.4800 ;
      RECT 0.4650 0.9000 0.5550 1.1750 ;
      RECT 0.0750 0.8100 0.5550 0.9000 ;
      RECT 0.0950 1.5700 0.2650 1.8250 ;
  END
END BUF_X1P4B_A12TH

MACRO BUF_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4300 0.3200 0.6000 0.7350 ;
        RECT 0.9500 0.3200 1.1200 0.7350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.4500 ;
        RECT 0.7300 1.4500 1.1500 1.5500 ;
        RECT 0.7250 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.5500 0.8200 1.9150 ;
        RECT 0.7250 0.4900 0.8250 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3500 1.3950 ;
    END
    ANTENNAGATEAREA 0.0402 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4700 1.7000 0.5600 2.0800 ;
        RECT 0.9900 1.7000 1.0800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4600 1.2550 0.9300 1.3450 ;
      RECT 0.1350 1.4850 0.5500 1.5750 ;
      RECT 0.4600 1.3450 0.5500 1.4850 ;
      RECT 0.4600 0.9200 0.5500 1.2550 ;
      RECT 0.1350 0.8300 0.5500 0.9200 ;
      RECT 0.1350 1.5750 0.2250 1.8900 ;
      RECT 0.1350 0.7100 0.2250 0.8300 ;
  END
END BUF_X1P4M_A12TH

MACRO BUF_X1P7B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4600 0.3200 0.5500 0.6100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4600 1.6750 0.5500 2.0800 ;
        RECT 0.9800 1.6750 1.0700 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.0100 0.3500 1.3700 ;
    END
    ANTENNAGATEAREA 0.0405 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.7200 1.2500 1.1500 1.3500 ;
        RECT 0.7150 0.8500 1.1500 0.9500 ;
        RECT 0.7200 1.3500 0.8100 1.7700 ;
        RECT 0.7150 0.5200 0.8150 0.8500 ;
    END
    ANTENNADIFFAREA 0.31085 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0700 0.9300 1.1600 ;
      RECT 0.1250 1.4800 0.5500 1.5700 ;
      RECT 0.4600 1.1600 0.5500 1.4800 ;
      RECT 0.4600 0.9000 0.5500 1.0700 ;
      RECT 0.0650 0.8100 0.5500 0.9000 ;
      RECT 0.1250 1.5700 0.2150 1.6900 ;
  END
END BUF_X1P7B_A12TH

MACRO BUF_X1P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4800 0.3200 0.5700 0.7300 ;
        RECT 1.0000 0.3200 1.0900 0.7300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3700 1.3600 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.7400 1.2500 1.1500 1.3500 ;
        RECT 0.7400 0.8500 1.1500 0.9500 ;
        RECT 0.7400 1.3500 0.8300 1.7150 ;
        RECT 0.7400 0.4900 0.8300 0.8500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4800 1.6600 0.5700 2.0800 ;
        RECT 1.0000 1.6250 1.0900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5200 1.0600 0.9400 1.1500 ;
      RECT 0.0650 1.4800 0.6100 1.5700 ;
      RECT 0.5200 1.1500 0.6100 1.4800 ;
      RECT 0.5200 0.9200 0.6100 1.0600 ;
      RECT 0.1250 0.8300 0.6100 0.9200 ;
      RECT 0.1250 0.5300 0.2150 0.8300 ;
  END
END BUF_X1P7M_A12TH

MACRO BUF_X2B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.4950 ;
        RECT 0.9900 0.3200 1.0800 0.4950 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4700 1.7700 0.5600 2.0800 ;
        RECT 0.9900 1.7700 1.0800 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7500 1.1500 1.2500 ;
        RECT 0.7300 1.2500 1.1500 1.3500 ;
        RECT 0.7250 0.6500 1.1500 0.7500 ;
        RECT 0.7300 1.3500 0.8200 1.7200 ;
        RECT 0.7250 0.5300 0.8250 0.6500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8100 0.3500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4800 1.0400 0.9400 1.1400 ;
      RECT 0.1350 1.2900 0.5700 1.3800 ;
      RECT 0.4800 1.1400 0.5700 1.2900 ;
      RECT 0.4800 0.7200 0.5700 1.0400 ;
      RECT 0.1350 0.6300 0.5700 0.7200 ;
      RECT 0.1350 1.3800 0.2250 1.7200 ;
      RECT 0.1350 0.5000 0.2250 0.6300 ;
  END
END BUF_X2B_A12TH

MACRO BUF_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.6300 ;
        RECT 0.9900 0.3200 1.0800 0.6300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.7300 1.2500 1.1500 1.3500 ;
        RECT 0.7250 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.3500 0.8200 1.7200 ;
        RECT 0.7250 0.4850 0.8250 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.4700 1.7700 0.5600 2.0800 ;
        RECT 0.9900 1.7700 1.0800 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0000 0.3600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4700 1.0600 0.9300 1.1500 ;
      RECT 0.1350 1.4800 0.5600 1.5700 ;
      RECT 0.4700 1.1500 0.5600 1.4800 ;
      RECT 0.4700 0.9050 0.5600 1.0600 ;
      RECT 0.1350 0.8150 0.5600 0.9050 ;
      RECT 0.1350 1.5700 0.2250 1.6900 ;
      RECT 0.1350 0.4950 0.2250 0.8150 ;
  END
END BUF_X2M_A12TH

MACRO BUF_X2P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4350 0.3200 0.5250 0.7350 ;
        RECT 0.9550 0.3200 1.0450 0.7550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.4350 1.6750 0.5250 2.0800 ;
        RECT 0.9550 1.6750 1.0450 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.3700 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.4500 ;
        RECT 0.6950 1.4500 1.3050 1.5500 ;
        RECT 0.6900 0.8500 1.1500 0.9500 ;
        RECT 0.6950 1.5500 0.7850 1.8800 ;
        RECT 1.2150 1.5500 1.3050 1.8800 ;
        RECT 0.6900 0.4850 0.7900 0.8500 ;
    END
    ANTENNADIFFAREA 0.399 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.4700 1.0600 0.9600 1.1500 ;
      RECT 0.0950 0.5900 0.2650 0.8250 ;
      RECT 0.1350 1.5700 0.2250 1.9100 ;
      RECT 0.1350 1.4800 0.5600 1.5700 ;
      RECT 0.4700 1.1500 0.5600 1.4800 ;
      RECT 0.4700 0.9150 0.5600 1.0600 ;
      RECT 0.0950 0.8250 0.5600 0.9150 ;
  END
END BUF_X2P5B_A12TH

MACRO BUF_X2P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4300 0.3200 0.5200 0.7250 ;
        RECT 0.9500 0.3200 1.0400 0.7250 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0681 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.2500 ;
        RECT 0.6900 1.2500 1.3500 1.3500 ;
        RECT 0.6850 0.8500 1.3500 0.9500 ;
        RECT 0.6900 1.3500 0.7800 1.7150 ;
        RECT 1.2100 1.3500 1.3000 1.7150 ;
        RECT 0.6850 0.4850 0.7850 0.8500 ;
        RECT 1.2100 0.4850 1.3000 0.8500 ;
    END
    ANTENNADIFFAREA 0.51 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3900 1.6800 0.5600 2.0800 ;
        RECT 0.9500 1.6200 1.0400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0600 1.0650 1.1500 ;
      RECT 0.0950 1.5700 0.1850 1.9100 ;
      RECT 0.0950 0.4850 0.1850 0.8250 ;
      RECT 0.0950 1.4800 0.5500 1.5700 ;
      RECT 0.4600 1.1500 0.5500 1.4800 ;
      RECT 0.4600 0.9150 0.5500 1.0600 ;
      RECT 0.0950 0.8250 0.5500 0.9150 ;
  END
END BUF_X2P5M_A12TH

MACRO BUF_X3B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4300 0.3200 0.5200 0.6700 ;
        RECT 0.9500 0.3200 1.0400 0.6700 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.4300 1.7700 0.5200 2.0800 ;
        RECT 0.9500 1.7700 1.0400 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0050 0.3600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0684 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.2500 ;
        RECT 0.6900 1.2500 1.3500 1.3500 ;
        RECT 0.6850 0.8500 1.3500 0.9500 ;
        RECT 0.6900 1.3500 0.7800 1.7150 ;
        RECT 1.2100 1.3500 1.3500 1.7150 ;
        RECT 0.6850 0.4850 0.7850 0.8500 ;
        RECT 1.2100 0.4850 1.3500 0.8500 ;
    END
    ANTENNADIFFAREA 0.511875 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.4700 1.0600 1.0800 1.1500 ;
      RECT 0.0950 1.5700 0.1850 1.9100 ;
      RECT 0.0950 0.5050 0.1850 0.8250 ;
      RECT 0.0950 1.4800 0.5600 1.5700 ;
      RECT 0.4700 1.1500 0.5600 1.4800 ;
      RECT 0.4700 0.9150 0.5600 1.0600 ;
      RECT 0.0950 0.8250 0.5600 0.9150 ;
  END
END BUF_X3B_A12TH

MACRO BUF_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.4300 0.3200 0.5200 0.6300 ;
        RECT 0.9500 0.3200 1.0400 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.4300 1.7700 0.5200 2.0800 ;
        RECT 0.9500 1.7700 1.0400 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.2500 ;
        RECT 0.6900 1.2500 1.3500 1.3500 ;
        RECT 0.6850 0.8500 1.3500 0.9500 ;
        RECT 0.6900 1.3500 0.7800 1.7200 ;
        RECT 1.2100 1.3500 1.3500 1.7200 ;
        RECT 0.6850 0.4850 0.7850 0.8500 ;
        RECT 1.2100 0.4850 1.3500 0.8500 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0801 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4700 1.0600 1.0700 1.1500 ;
      RECT 0.0950 1.5700 0.1850 1.9100 ;
      RECT 0.0950 0.4950 0.1850 0.8250 ;
      RECT 0.0950 1.4800 0.5600 1.5700 ;
      RECT 0.4700 1.1500 0.5600 1.4800 ;
      RECT 0.4700 0.9150 0.5600 1.0600 ;
      RECT 0.0950 0.8250 0.5600 0.9150 ;
  END
END BUF_X3M_A12TH

MACRO BUF_X3P5B_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6400 ;
        RECT 0.8500 0.3200 1.0200 0.7550 ;
        RECT 1.3700 0.3200 1.5400 0.7550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3500 1.6800 0.4500 2.0800 ;
        RECT 0.8850 1.6550 0.9850 2.0800 ;
        RECT 1.4050 1.6550 1.5050 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9800 0.3500 1.3700 ;
    END
    ANTENNAGATEAREA 0.0801 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.2500 ;
        RECT 0.6300 1.2500 1.3500 1.3500 ;
        RECT 0.6300 0.8500 1.3500 0.9500 ;
        RECT 0.6300 1.3500 0.7200 1.7200 ;
        RECT 1.1500 1.3500 1.2400 1.7200 ;
        RECT 0.6300 0.4400 0.7200 0.8500 ;
        RECT 1.1500 0.4400 1.2400 0.8500 ;
    END
    ANTENNADIFFAREA 0.478 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.4500 1.0600 1.0700 1.1500 ;
      RECT 0.0950 1.5900 0.1850 1.9300 ;
      RECT 0.0950 0.4400 0.1850 0.7700 ;
      RECT 0.0950 1.5000 0.5400 1.5900 ;
      RECT 0.4500 1.1500 0.5400 1.5000 ;
      RECT 0.4500 0.8600 0.5400 1.0600 ;
      RECT 0.0950 0.7700 0.5400 0.8600 ;
  END
END BUF_X3P5B_A12TH

MACRO BUF_X3P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6900 ;
        RECT 0.8900 0.3200 0.9800 0.6950 ;
        RECT 1.4100 0.3200 1.5000 0.6950 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3550 1.6800 0.4450 2.0800 ;
        RECT 0.8900 1.6550 0.9800 2.0800 ;
        RECT 1.4100 1.6550 1.5000 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.4500 ;
        RECT 0.6300 1.4500 1.3500 1.5500 ;
        RECT 0.6300 0.8500 1.3500 0.9500 ;
        RECT 0.6300 1.5500 0.7200 1.8800 ;
        RECT 1.1500 1.5500 1.2400 1.8800 ;
        RECT 0.6300 0.4600 0.7200 0.8500 ;
        RECT 1.1500 0.4600 1.2400 0.8500 ;
    END
    ANTENNADIFFAREA 0.568 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3600 1.3700 ;
    END
    ANTENNAGATEAREA 0.0939 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4500 1.0600 1.0700 1.1500 ;
      RECT 0.0950 1.5900 0.1850 1.9300 ;
      RECT 0.0950 0.4600 0.1850 0.8100 ;
      RECT 0.0950 1.5000 0.5400 1.5900 ;
      RECT 0.4500 1.1500 0.5400 1.5000 ;
      RECT 0.4500 0.9000 0.5400 1.0600 ;
      RECT 0.0950 0.8100 0.5400 0.9000 ;
  END
END BUF_X3P5M_A12TH

MACRO BUFH_X0P8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3700 0.3200 0.4600 0.4700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6300 0.4850 0.7500 1.7200 ;
    END
    ANTENNADIFFAREA 0.2184 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8000 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3650 1.6400 0.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.3000 0.5350 1.3900 ;
      RECT 0.4450 0.6800 0.5350 1.3000 ;
      RECT 0.0750 0.5900 0.5350 0.6800 ;
      RECT 0.0750 1.3900 0.1750 1.7300 ;
      RECT 0.0750 0.4900 0.1750 0.5900 ;
  END
END BUFH_X0P8M_A12TH

MACRO BUFH_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.6600 ;
        RECT 0.6450 0.3200 0.7350 0.6600 ;
        RECT 1.1650 0.3200 1.2550 0.6600 ;
        RECT 1.6900 0.3200 1.7800 0.6600 ;
        RECT 2.2200 0.3200 2.3100 0.6600 ;
        RECT 2.7400 0.3200 2.8300 0.6600 ;
        RECT 3.2600 0.3200 3.3500 0.6600 ;
        RECT 3.7800 0.3200 3.8700 0.6600 ;
        RECT 4.3000 0.3200 4.3900 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.1250 1.7700 0.2150 2.0800 ;
        RECT 0.6450 1.7700 0.7350 2.0800 ;
        RECT 1.1650 1.7700 1.2550 2.0800 ;
        RECT 1.6900 1.7700 1.7800 2.0800 ;
        RECT 2.2200 1.7700 2.3100 2.0800 ;
        RECT 2.7400 1.7700 2.8300 2.0800 ;
        RECT 3.2600 1.7700 3.3500 2.0800 ;
        RECT 3.7800 1.7700 3.8700 2.0800 ;
        RECT 4.3000 1.7700 4.3900 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4200 0.9800 4.5800 1.4200 ;
        RECT 1.9600 1.4200 4.6500 1.5800 ;
        RECT 1.9600 0.8200 4.6500 0.9800 ;
        RECT 1.9600 1.5800 2.0500 1.8500 ;
        RECT 2.4800 1.5800 2.5700 1.8500 ;
        RECT 3.0000 1.5800 3.0900 1.8500 ;
        RECT 3.5200 1.5800 3.6100 1.8500 ;
        RECT 4.0400 1.5800 4.1300 1.8500 ;
        RECT 4.5600 1.5800 4.6500 1.8500 ;
        RECT 1.9600 0.5150 2.0500 0.8200 ;
        RECT 2.4800 0.5150 2.5700 0.8200 ;
        RECT 3.0000 0.5150 3.0900 0.8200 ;
        RECT 3.5200 0.5150 3.6100 0.8200 ;
        RECT 4.0400 0.5150 4.1300 0.8200 ;
        RECT 4.5600 0.5150 4.6500 0.8200 ;
    END
    ANTENNADIFFAREA 1.958125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0500 1.4500 1.1500 ;
    END
    ANTENNAGATEAREA 0.585 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.7000 1.0700 4.0550 1.1600 ;
      RECT 0.3850 1.3700 0.4750 1.7200 ;
      RECT 0.3850 0.4900 0.4750 0.8300 ;
      RECT 0.9050 1.3700 0.9950 1.7200 ;
      RECT 0.9050 0.4900 0.9950 0.8300 ;
      RECT 1.4250 1.3700 1.5150 1.7200 ;
      RECT 1.4250 0.4900 1.5150 0.8300 ;
      RECT 0.3850 1.2800 1.7900 1.3700 ;
      RECT 1.7000 1.1600 1.7900 1.2800 ;
      RECT 1.7000 0.9200 1.7900 1.0700 ;
      RECT 0.3850 0.8300 1.7900 0.9200 ;
  END
END BUFH_X11M_A12TH

MACRO BUFH_X13M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7200 ;
        RECT 0.6150 0.3200 0.7050 0.7200 ;
        RECT 1.1350 0.3200 1.2250 0.7200 ;
        RECT 1.6550 0.3200 1.7450 0.7200 ;
        RECT 2.1750 0.3200 2.2650 0.7200 ;
        RECT 2.7100 0.3200 2.8000 0.6600 ;
        RECT 3.2300 0.3200 3.3200 0.6600 ;
        RECT 3.7500 0.3200 3.8400 0.6600 ;
        RECT 4.2700 0.3200 4.3600 0.6600 ;
        RECT 4.7900 0.3200 4.8800 0.6600 ;
        RECT 5.3100 0.3200 5.4000 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 2.7100 1.7700 2.8000 2.0800 ;
        RECT 3.2300 1.7700 3.3200 2.0800 ;
        RECT 3.7500 1.7700 3.8400 2.0800 ;
        RECT 4.2700 1.7700 4.3600 2.0800 ;
        RECT 4.7900 1.7700 4.8800 2.0800 ;
        RECT 5.3100 1.7700 5.4000 2.0800 ;
        RECT 0.0900 1.6900 0.1800 2.0800 ;
        RECT 0.6150 1.6900 0.7050 2.0800 ;
        RECT 1.1350 1.6900 1.2250 2.0800 ;
        RECT 1.6550 1.6900 1.7450 2.0800 ;
        RECT 2.1800 1.6900 2.2700 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4100 0.9900 5.5900 1.4100 ;
        RECT 2.4500 1.4100 5.6600 1.5900 ;
        RECT 2.4500 0.8100 5.6600 0.9900 ;
        RECT 2.4500 1.5900 2.5400 1.8400 ;
        RECT 2.9700 1.5900 3.0600 1.8400 ;
        RECT 3.4900 1.5900 3.5800 1.8400 ;
        RECT 4.0100 1.5900 4.1000 1.8400 ;
        RECT 4.5300 1.5900 4.6200 1.8400 ;
        RECT 5.0500 1.5900 5.1400 1.8400 ;
        RECT 5.5700 1.5900 5.6600 1.8400 ;
        RECT 2.4500 0.5150 2.5400 0.8100 ;
        RECT 2.9700 0.5150 3.0600 0.8100 ;
        RECT 3.4900 0.5150 3.5800 0.8100 ;
        RECT 4.0100 0.5150 4.1000 0.8100 ;
        RECT 4.5300 0.5150 4.6200 0.8100 ;
        RECT 5.0500 0.5150 5.1400 0.8100 ;
        RECT 5.5700 0.5150 5.6600 0.8100 ;
    END
    ANTENNADIFFAREA 2.283125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 1.0500 1.8250 1.1500 ;
    END
    ANTENNAGATEAREA 0.7128 ;
  END A
  OBS
    LAYER M1 ;
      RECT 2.2200 1.0800 4.6900 1.1700 ;
      RECT 0.3550 1.3700 0.4450 1.7200 ;
      RECT 0.3550 0.4900 0.4450 0.8300 ;
      RECT 0.8750 1.3700 0.9650 1.7200 ;
      RECT 0.8750 0.4900 0.9650 0.8300 ;
      RECT 1.3950 1.3700 1.4850 1.7200 ;
      RECT 1.3950 0.4900 1.4850 0.8300 ;
      RECT 1.9150 1.3700 2.0050 1.7200 ;
      RECT 1.9150 0.4900 2.0050 0.8300 ;
      RECT 0.3550 1.2800 2.3100 1.3700 ;
      RECT 2.2200 1.1700 2.3100 1.2800 ;
      RECT 2.2200 0.9200 2.3100 1.0800 ;
      RECT 0.3550 0.8300 2.3100 0.9200 ;
  END
END BUFH_X13M_A12TH

MACRO BUFH_X16M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6600 ;
        RECT 0.8750 0.3200 0.9650 0.6600 ;
        RECT 1.3950 0.3200 1.4850 0.6600 ;
        RECT 1.9150 0.3200 2.0050 0.6600 ;
        RECT 2.4350 0.3200 2.5250 0.6600 ;
        RECT 2.9700 0.3200 3.0600 0.6600 ;
        RECT 3.4900 0.3200 3.5800 0.6600 ;
        RECT 4.0100 0.3200 4.1000 0.6600 ;
        RECT 4.5300 0.3200 4.6200 0.6600 ;
        RECT 5.0500 0.3200 5.1400 0.6600 ;
        RECT 5.5700 0.3200 5.6600 0.6600 ;
        RECT 6.0900 0.3200 6.1800 0.6600 ;
        RECT 6.6100 0.3200 6.7000 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
        RECT 1.9150 1.7700 2.0050 2.0800 ;
        RECT 2.4500 1.7700 2.5400 2.0800 ;
        RECT 2.9700 1.7700 3.0600 2.0800 ;
        RECT 3.4900 1.7700 3.5800 2.0800 ;
        RECT 4.0100 1.7700 4.1000 2.0800 ;
        RECT 4.5300 1.7700 4.6200 2.0800 ;
        RECT 5.0500 1.7700 5.1400 2.0800 ;
        RECT 5.5700 1.7700 5.6600 2.0800 ;
        RECT 6.0900 1.7700 6.1800 2.0800 ;
        RECT 6.6100 1.7700 6.7000 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.1900 1.0000 6.4400 1.3900 ;
        RECT 2.7100 1.3900 6.4400 1.6100 ;
        RECT 2.7100 0.7800 6.4400 1.0000 ;
        RECT 2.7100 1.6100 2.8000 1.8250 ;
        RECT 3.2300 1.6100 3.3200 1.8250 ;
        RECT 3.7500 1.6100 3.8400 1.8250 ;
        RECT 4.2700 1.6100 4.3600 1.8250 ;
        RECT 4.7900 1.6100 4.8800 1.8250 ;
        RECT 5.3100 1.6100 5.4000 1.8250 ;
        RECT 5.8300 1.6100 5.9200 1.8250 ;
        RECT 6.3500 1.6100 6.4400 1.8250 ;
        RECT 2.7100 0.5150 2.8000 0.7800 ;
        RECT 3.2300 0.5150 3.3200 0.7800 ;
        RECT 3.7500 0.5150 3.8400 0.7800 ;
        RECT 4.2700 0.5150 4.3600 0.7800 ;
        RECT 4.7900 0.5150 4.8800 0.7800 ;
        RECT 5.3100 0.5150 5.4000 0.7800 ;
        RECT 5.8300 0.5150 5.9200 0.7800 ;
        RECT 6.3500 0.5150 6.4400 0.7800 ;
    END
    ANTENNADIFFAREA 2.6 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3000 1.0500 2.0750 1.1500 ;
    END
    ANTENNAGATEAREA 0.8775 ;
  END A
  OBS
    LAYER M1 ;
      RECT 2.4800 1.1100 5.6150 1.2000 ;
      RECT 0.0950 1.3700 0.1850 1.7200 ;
      RECT 0.0950 0.4900 0.1850 0.8300 ;
      RECT 0.6150 1.3700 0.7050 1.7200 ;
      RECT 0.6150 0.4900 0.7050 0.8300 ;
      RECT 1.1350 1.3700 1.2250 1.7200 ;
      RECT 1.1350 0.4900 1.2250 0.8300 ;
      RECT 1.6550 1.3700 1.7450 1.7200 ;
      RECT 1.6550 0.4900 1.7450 0.8300 ;
      RECT 2.1750 1.3700 2.2650 1.7200 ;
      RECT 2.1750 0.4900 2.2650 0.8300 ;
      RECT 0.0950 1.2800 2.5700 1.3700 ;
      RECT 2.4800 1.2000 2.5700 1.2800 ;
      RECT 2.4800 0.9200 2.5700 1.1100 ;
      RECT 0.0950 0.8300 2.5700 0.9200 ;
  END
END BUFH_X16M_A12TH

MACRO BUFH_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.7900 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8950 0.7500 1.4750 ;
        RECT 0.6300 1.4750 0.7500 1.8850 ;
        RECT 0.6300 0.4850 0.7500 0.8950 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3650 1.7700 0.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.3000 0.5350 1.3900 ;
      RECT 0.4450 0.6400 0.5350 1.3000 ;
      RECT 0.0750 0.5500 0.5350 0.6400 ;
      RECT 0.0550 1.3900 0.1750 1.7300 ;
      RECT 0.0750 0.4300 0.1750 0.5500 ;
  END
END BUFH_X1M_A12TH

MACRO BUFH_X1P2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7350 ;
        RECT 0.9900 0.3200 1.0800 0.7300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.4500 ;
        RECT 0.7300 1.4500 1.1500 1.5500 ;
        RECT 0.7300 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.5500 0.8200 1.8800 ;
        RECT 0.7300 0.5100 0.8200 0.8500 ;
    END
    ANTENNADIFFAREA 0.193 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3950 1.6700 0.4850 2.0800 ;
        RECT 0.9500 1.6550 1.1200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0600 0.9300 1.1500 ;
      RECT 0.1350 1.4800 0.5500 1.5700 ;
      RECT 0.4600 1.1500 0.5500 1.4800 ;
      RECT 0.4600 0.9150 0.5500 1.0600 ;
      RECT 0.1350 0.8250 0.5500 0.9150 ;
      RECT 0.1350 1.5700 0.2250 1.9100 ;
      RECT 0.1350 0.4800 0.2250 0.8250 ;
  END
END BUFH_X1P2M_A12TH

MACRO BUFH_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.4050 0.3200 0.4950 0.7350 ;
        RECT 0.9450 0.3200 1.1150 0.7400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3650 1.6900 0.5350 2.0800 ;
        RECT 0.9850 1.5250 1.0750 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9450 1.1500 1.2500 ;
        RECT 0.7250 1.2500 1.1500 1.3500 ;
        RECT 0.7250 0.8550 1.1500 0.9450 ;
        RECT 0.7250 1.3500 0.8150 1.7200 ;
        RECT 0.7250 0.5150 0.8150 0.8550 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0650 0.9250 1.1550 ;
      RECT 0.1450 1.4800 0.5500 1.5700 ;
      RECT 0.4600 1.1550 0.5500 1.4800 ;
      RECT 0.4600 0.9150 0.5500 1.0650 ;
      RECT 0.1450 0.8250 0.5500 0.9150 ;
      RECT 0.1450 1.5700 0.2350 1.9100 ;
      RECT 0.1450 0.4850 0.2350 0.8250 ;
  END
END BUFH_X1P4M_A12TH

MACRO BUFH_X1P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.3950 0.3200 0.4850 0.6900 ;
        RECT 0.9900 0.3200 1.0800 0.7550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3950 1.7300 0.4850 2.0800 ;
        RECT 0.9900 1.6250 1.0800 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0933 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9500 1.1500 1.2500 ;
        RECT 0.7300 1.2500 1.1500 1.3500 ;
        RECT 0.7300 0.8500 1.1500 0.9500 ;
        RECT 0.7300 1.3500 0.8200 1.7200 ;
        RECT 0.7300 0.5150 0.8200 0.8500 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0650 0.9300 1.1550 ;
      RECT 0.1350 1.4800 0.5500 1.5700 ;
      RECT 0.4600 1.1550 0.5500 1.4800 ;
      RECT 0.4600 0.9150 0.5500 1.0650 ;
      RECT 0.1350 0.8250 0.5500 0.9150 ;
      RECT 0.1350 1.5700 0.2250 1.9100 ;
      RECT 0.1350 0.5050 0.2250 0.8250 ;
  END
END BUFH_X1P7M_A12TH

MACRO BUFH_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.9550 ;
        RECT 0.6900 0.3200 0.7800 0.6600 ;
        RECT 1.2100 0.3200 1.3000 0.6600 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1116 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.2500 ;
        RECT 0.9500 1.2500 1.3500 1.3500 ;
        RECT 0.9500 0.8500 1.3500 0.9500 ;
        RECT 0.9500 1.3500 1.0400 1.7200 ;
        RECT 0.9500 0.5150 1.0400 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6900 1.7700 0.7800 2.0800 ;
        RECT 1.2100 1.7700 1.3000 2.0800 ;
        RECT 0.0950 1.3800 0.1850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7000 1.0650 1.1300 1.1550 ;
      RECT 0.3550 1.2800 0.7900 1.3700 ;
      RECT 0.7000 1.1550 0.7900 1.2800 ;
      RECT 0.7000 0.9200 0.7900 1.0650 ;
      RECT 0.3550 0.8300 0.7900 0.9200 ;
      RECT 0.3550 1.3700 0.4450 1.7200 ;
      RECT 0.3550 0.4900 0.4450 0.8300 ;
  END
END BUFH_X2M_A12TH

MACRO BUFH_X2P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.8650 ;
        RECT 0.5750 0.3200 0.7450 0.7400 ;
        RECT 1.1500 0.3200 1.2400 0.7550 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1500 1.6200 1.2400 2.0800 ;
        RECT 0.0950 1.5100 0.1850 2.0800 ;
        RECT 0.6150 1.5100 0.7050 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.2500 ;
        RECT 0.8900 1.2500 1.5500 1.3500 ;
        RECT 0.8900 0.8500 1.5500 0.9500 ;
        RECT 0.8900 1.3500 0.9800 1.7200 ;
        RECT 1.4100 1.3500 1.5500 1.7200 ;
        RECT 0.8900 0.5150 0.9800 0.8500 ;
        RECT 1.4100 0.5150 1.5500 0.8500 ;
    END
    ANTENNADIFFAREA 0.51 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.6900 1.0650 1.2500 1.1550 ;
      RECT 0.3550 1.3700 0.4450 1.7200 ;
      RECT 0.3550 0.4900 0.4450 0.8300 ;
      RECT 0.3550 1.2800 0.7800 1.3700 ;
      RECT 0.6900 1.1550 0.7800 1.2800 ;
      RECT 0.6900 0.9200 0.7800 1.0650 ;
      RECT 0.3550 0.8300 0.7800 0.9200 ;
  END
END BUFH_X2P5M_A12TH

MACRO BUFH_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7750 ;
        RECT 0.6150 0.3200 0.7050 0.7350 ;
        RECT 1.1500 0.3200 1.2400 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1500 1.7700 1.2400 2.0800 ;
        RECT 0.0950 1.6200 0.1850 2.0800 ;
        RECT 0.6150 1.6200 0.7050 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5500 1.2500 ;
        RECT 0.8900 1.2500 1.5500 1.3500 ;
        RECT 0.8900 0.8500 1.5500 0.9500 ;
        RECT 0.8900 1.3500 0.9800 1.7200 ;
        RECT 1.4100 1.3500 1.5500 1.7250 ;
        RECT 0.8900 0.5150 0.9800 0.8500 ;
        RECT 1.4100 0.5150 1.5500 0.8500 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1632 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.6900 1.0650 1.2450 1.1550 ;
      RECT 0.3550 1.3700 0.4450 1.7050 ;
      RECT 0.3550 0.5000 0.4450 0.8300 ;
      RECT 0.3550 1.2800 0.7800 1.3700 ;
      RECT 0.6900 1.1550 0.7800 1.2800 ;
      RECT 0.6900 0.9200 0.7800 1.0650 ;
      RECT 0.3550 0.8300 0.7800 0.9200 ;
  END
END BUFH_X3M_A12TH

MACRO BUFH_X3P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6750 ;
        RECT 0.6150 0.3200 0.7050 0.7300 ;
        RECT 1.1500 0.3200 1.2400 0.7500 ;
        RECT 1.6700 0.3200 1.7600 0.7500 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1200 1.0500 0.5400 1.1500 ;
    END
    ANTENNAGATEAREA 0.1908 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.0950 1.7500 0.1850 2.0800 ;
        RECT 0.6150 1.6550 0.7050 2.0800 ;
        RECT 1.1500 1.6550 1.2400 2.0800 ;
        RECT 1.6700 1.6550 1.7600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.2500 ;
        RECT 0.8900 1.2500 1.7500 1.3500 ;
        RECT 0.8900 0.8500 1.7500 0.9500 ;
        RECT 0.8900 1.3500 0.9800 1.7200 ;
        RECT 1.4100 1.3500 1.5000 1.7250 ;
        RECT 0.8900 0.5150 0.9800 0.8500 ;
        RECT 1.4100 0.5150 1.5000 0.8500 ;
    END
    ANTENNADIFFAREA 0.568 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.6900 1.0650 1.4550 1.1550 ;
      RECT 0.3550 1.3700 0.4450 1.7200 ;
      RECT 0.3550 0.4900 0.4450 0.8300 ;
      RECT 0.3550 1.2800 0.7800 1.3700 ;
      RECT 0.6900 1.1550 0.7800 1.2800 ;
      RECT 0.6900 0.9200 0.7800 1.0650 ;
      RECT 0.3550 0.8300 0.7800 0.9200 ;
  END
END BUFH_X3P5M_A12TH

MACRO BUFH_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.3450 0.3200 0.5150 0.7100 ;
        RECT 0.8650 0.3200 1.0350 0.7100 ;
        RECT 1.4400 0.3200 1.5300 0.6600 ;
        RECT 1.9600 0.3200 2.0500 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.4400 1.7700 1.5300 2.0800 ;
        RECT 1.9600 1.7700 2.0500 2.0800 ;
        RECT 0.3850 1.5500 0.4750 2.0800 ;
        RECT 0.9050 1.5500 0.9950 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9500 1.9500 1.2500 ;
        RECT 1.1800 1.2500 1.9500 1.3500 ;
        RECT 1.1800 0.8500 1.9500 0.9500 ;
        RECT 1.1800 1.3500 1.2700 1.7250 ;
        RECT 1.7000 1.3500 1.7900 1.7250 ;
        RECT 1.1800 0.5150 1.2700 0.8500 ;
        RECT 1.7000 0.5150 1.7900 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.0500 0.7550 1.1500 ;
    END
    ANTENNAGATEAREA 0.2223 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.9000 1.0650 1.7000 1.1550 ;
      RECT 0.1250 1.3700 0.2150 1.7200 ;
      RECT 0.1250 0.4900 0.2150 0.8300 ;
      RECT 0.6450 1.3700 0.7350 1.7200 ;
      RECT 0.6450 0.4900 0.7350 0.8300 ;
      RECT 0.1250 1.2800 0.9900 1.3700 ;
      RECT 0.9000 1.1550 0.9900 1.2800 ;
      RECT 0.9000 0.9200 0.9900 1.0650 ;
      RECT 0.1250 0.8300 0.9900 0.9200 ;
  END
END BUFH_X4M_A12TH

MACRO BUFH_X5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3800 0.3200 0.4700 0.7050 ;
        RECT 0.9000 0.3200 0.9900 0.7050 ;
        RECT 1.4350 0.3200 1.5250 0.6600 ;
        RECT 1.9550 0.3200 2.0450 0.6600 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0500 0.7500 1.1500 ;
    END
    ANTENNAGATEAREA 0.2736 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.2500 ;
        RECT 1.1750 1.2500 2.3500 1.3500 ;
        RECT 1.1750 0.8500 2.3500 0.9500 ;
        RECT 1.1750 1.3500 1.2650 1.7200 ;
        RECT 1.6950 1.3500 1.7850 1.7200 ;
        RECT 2.2150 1.3500 2.3050 1.7200 ;
        RECT 1.1750 0.5150 1.2650 0.8500 ;
        RECT 1.6950 0.5150 1.7850 0.8500 ;
        RECT 2.2150 0.5150 2.3050 0.8500 ;
    END
    ANTENNADIFFAREA 0.934375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 1.4350 1.7700 1.5250 2.0800 ;
        RECT 1.9550 1.7700 2.0450 2.0800 ;
        RECT 0.3800 1.7100 0.4700 2.0800 ;
        RECT 0.9050 1.7100 0.9950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.9000 1.0650 2.0500 1.1550 ;
      RECT 0.1200 1.3700 0.2100 1.7200 ;
      RECT 0.1200 0.4900 0.2100 0.8300 ;
      RECT 0.6400 1.3700 0.7300 1.7200 ;
      RECT 0.6400 0.4900 0.7300 0.8300 ;
      RECT 0.1200 1.2800 0.9900 1.3700 ;
      RECT 0.9000 1.1550 0.9900 1.2800 ;
      RECT 0.9000 0.9200 0.9900 1.0650 ;
      RECT 0.1200 0.8300 0.9900 0.9200 ;
  END
END BUFH_X5M_A12TH

MACRO BUFH_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.7700 ;
        RECT 0.6450 0.3200 0.7350 0.7400 ;
        RECT 1.1650 0.3200 1.2550 0.7400 ;
        RECT 1.7000 0.3200 1.7900 0.6600 ;
        RECT 2.2200 0.3200 2.3100 0.6600 ;
        RECT 2.7400 0.3200 2.8300 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 1.7000 1.7700 1.7900 2.0800 ;
        RECT 2.2200 1.7700 2.3100 2.0800 ;
        RECT 2.7400 1.7700 2.8300 2.0800 ;
        RECT 0.1250 1.6250 0.2150 2.0800 ;
        RECT 0.6450 1.6250 0.7350 2.0800 ;
        RECT 1.1700 1.6250 1.2600 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.0500 1.0050 1.1500 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9500 2.7500 1.2500 ;
        RECT 1.4400 1.2500 2.7500 1.3500 ;
        RECT 1.4400 0.8500 2.7500 0.9500 ;
        RECT 1.4400 1.3500 1.5300 1.7200 ;
        RECT 1.9600 1.3500 2.0500 1.7200 ;
        RECT 2.4800 1.3500 2.5700 1.7200 ;
        RECT 1.4400 0.5150 1.5300 0.8500 ;
        RECT 1.9600 0.5150 2.0500 0.8500 ;
        RECT 2.4800 0.5150 2.5700 0.8500 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.2400 1.0650 2.3750 1.1550 ;
      RECT 0.3850 1.3700 0.4750 1.7200 ;
      RECT 0.3850 0.4900 0.4750 0.8300 ;
      RECT 0.9050 1.3700 0.9950 1.7200 ;
      RECT 0.9050 0.4900 0.9950 0.8300 ;
      RECT 0.3850 1.2800 1.3300 1.3700 ;
      RECT 1.2400 1.1550 1.3300 1.2800 ;
      RECT 1.2400 0.9200 1.3300 1.0650 ;
      RECT 0.3850 0.8300 1.3300 0.9200 ;
  END
END BUFH_X6M_A12TH

MACRO BUFH_X7P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.3850 0.3200 0.4750 0.7400 ;
        RECT 0.9050 0.3200 0.9950 0.7400 ;
        RECT 1.4250 0.3200 1.5150 0.7400 ;
        RECT 1.9600 0.3200 2.0500 0.7000 ;
        RECT 2.4800 0.3200 2.5700 0.7000 ;
        RECT 3.0000 0.3200 3.0900 0.7000 ;
        RECT 3.5200 0.3200 3.6100 0.7000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 1.9600 1.7150 2.0500 2.0800 ;
        RECT 2.4800 1.7150 2.5700 2.0800 ;
        RECT 3.0000 1.7150 3.0900 2.0800 ;
        RECT 3.5200 1.7150 3.6100 2.0800 ;
        RECT 0.3850 1.6450 0.4750 2.0800 ;
        RECT 0.9050 1.6450 0.9950 2.0800 ;
        RECT 1.4250 1.6450 1.5150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2400 0.9600 3.3600 1.2400 ;
        RECT 1.7000 1.2400 3.3600 1.3600 ;
        RECT 1.7000 0.8400 3.3600 0.9600 ;
        RECT 1.7000 1.3600 1.7900 1.7250 ;
        RECT 2.2200 1.3600 2.3100 1.7250 ;
        RECT 2.7400 1.3600 2.8300 1.7250 ;
        RECT 3.2600 1.3600 3.3600 1.7250 ;
        RECT 1.7000 0.5150 1.7900 0.8400 ;
        RECT 2.2200 0.5150 2.3100 0.8400 ;
        RECT 2.7400 0.5150 2.8300 0.8400 ;
        RECT 3.2600 0.5150 3.3600 0.8400 ;
    END
    ANTENNADIFFAREA 1.224 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3800 1.0500 1.1900 1.1500 ;
    END
    ANTENNAGATEAREA 0.42 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.4600 1.0600 2.8400 1.1500 ;
      RECT 0.1250 1.3700 0.2150 1.7200 ;
      RECT 0.1250 0.4900 0.2150 0.8300 ;
      RECT 0.6450 1.3700 0.7350 1.7200 ;
      RECT 0.6450 0.4900 0.7350 0.8300 ;
      RECT 1.1650 1.3700 1.2550 1.7200 ;
      RECT 1.1650 0.4900 1.2550 0.8300 ;
      RECT 0.1250 1.2800 1.5500 1.3700 ;
      RECT 1.4600 1.1500 1.5500 1.2800 ;
      RECT 1.4600 0.9200 1.5500 1.0600 ;
      RECT 0.1250 0.8300 1.5500 0.9200 ;
  END
END BUFH_X7P5M_A12TH

MACRO BUFH_X9M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.3850 0.3200 0.4750 0.6600 ;
        RECT 0.9050 0.3200 0.9950 0.6600 ;
        RECT 1.4250 0.3200 1.5150 0.6600 ;
        RECT 1.9600 0.3200 2.0500 0.6600 ;
        RECT 2.4800 0.3200 2.5700 0.6600 ;
        RECT 3.0000 0.3200 3.0900 0.6600 ;
        RECT 3.5200 0.3200 3.6100 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.3850 1.7700 0.4750 2.0800 ;
        RECT 0.9050 1.7700 0.9950 2.0800 ;
        RECT 1.4300 1.7700 1.5200 2.0800 ;
        RECT 1.9600 1.7700 2.0500 2.0800 ;
        RECT 2.4800 1.7700 2.5700 2.0800 ;
        RECT 3.0000 1.7700 3.0900 2.0800 ;
        RECT 3.5200 1.7700 3.6100 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.0500 1.2100 1.1500 ;
    END
    ANTENNAGATEAREA 0.4875 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6350 0.9650 3.7650 1.2350 ;
        RECT 1.7000 1.2350 3.8700 1.3650 ;
        RECT 1.7000 0.8350 3.8700 0.9650 ;
        RECT 1.7000 1.3650 1.7900 1.7200 ;
        RECT 2.2200 1.3650 2.3100 1.7200 ;
        RECT 2.7400 1.3650 2.8300 1.7200 ;
        RECT 3.2600 1.3650 3.3500 1.7200 ;
        RECT 3.7800 1.3650 3.8700 1.7200 ;
        RECT 1.7000 0.5150 1.7900 0.8350 ;
        RECT 2.2200 0.5150 2.3100 0.8350 ;
        RECT 2.7400 0.5150 2.8300 0.8350 ;
        RECT 3.2600 0.5150 3.3500 0.8350 ;
        RECT 3.7800 0.5150 3.8700 0.8350 ;
    END
    ANTENNADIFFAREA 1.616225 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.4800 1.0550 3.3250 1.1450 ;
      RECT 0.6450 1.3700 0.7350 1.7200 ;
      RECT 0.6450 0.4900 0.7350 0.8300 ;
      RECT 1.1650 1.3700 1.2550 1.7200 ;
      RECT 1.1650 0.4900 1.2550 0.8300 ;
      RECT 0.1250 1.2800 1.5700 1.3700 ;
      RECT 1.4800 1.1450 1.5700 1.2800 ;
      RECT 1.4800 0.9200 1.5700 1.0550 ;
      RECT 0.1250 0.8300 1.5700 0.9200 ;
      RECT 0.1250 1.3700 0.2150 1.7200 ;
      RECT 0.1250 0.4900 0.2150 0.8300 ;
  END
END BUFH_X9M_A12TH

MACRO BUFZ_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.1100 0.3200 0.2000 0.6900 ;
        RECT 0.5900 0.3200 0.7600 0.5650 ;
        RECT 1.1250 0.3200 1.2950 0.3950 ;
        RECT 2.7600 0.3200 2.8500 0.6450 ;
        RECT 3.2800 0.3200 3.3700 0.6450 ;
        RECT 3.8000 0.3200 3.8900 0.6550 ;
        RECT 4.3500 0.3200 4.4400 0.6300 ;
        RECT 4.8300 0.3200 5.0000 0.5700 ;
        RECT 5.3500 0.3200 5.5200 0.5700 ;
        RECT 5.8700 0.3200 6.0400 0.5700 ;
        RECT 6.3900 0.3200 6.5600 0.5700 ;
        RECT 6.9100 0.3200 7.0800 0.5700 ;
        RECT 7.4300 0.3200 7.6000 0.5700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6700 1.4200 7.3600 1.5800 ;
        RECT 4.6700 1.5800 4.7600 1.8500 ;
        RECT 5.1900 1.5800 5.2800 1.8500 ;
        RECT 5.7100 1.5800 5.8000 1.8500 ;
        RECT 6.2300 1.5800 6.3200 1.8500 ;
        RECT 6.7500 1.5800 6.8400 1.8500 ;
        RECT 7.2700 1.5800 7.3600 1.8500 ;
        RECT 7.0200 0.8400 7.1800 1.4200 ;
        RECT 4.6100 0.6800 7.3000 0.8400 ;
        RECT 4.6100 0.4100 4.7000 0.6800 ;
        RECT 5.1300 0.4100 5.2200 0.6800 ;
        RECT 5.6500 0.4100 5.7400 0.6800 ;
        RECT 6.1700 0.4100 6.2600 0.6800 ;
        RECT 6.6900 0.4100 6.7800 0.6800 ;
        RECT 7.2100 0.4100 7.3000 0.6800 ;
    END
    ANTENNADIFFAREA 1.758 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7300 1.0500 3.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.4734 ;
  END A

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3400 1.0500 0.7500 1.1500 ;
        RECT 0.6500 0.8000 0.7500 1.0500 ;
        RECT 0.6500 0.7000 1.3750 0.8000 ;
        RECT 1.2850 0.8000 1.3750 1.0200 ;
    END
    ANTENNAGATEAREA 0.3687 ;
  END OE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 4.4100 1.7700 4.5000 2.0800 ;
        RECT 4.9300 1.7700 5.0200 2.0800 ;
        RECT 5.4500 1.7700 5.5400 2.0800 ;
        RECT 5.9700 1.7700 6.0600 2.0800 ;
        RECT 6.4900 1.7700 6.5800 2.0800 ;
        RECT 7.0100 1.7700 7.1000 2.0800 ;
        RECT 7.5300 1.7700 7.6200 2.0800 ;
        RECT 0.1100 1.7100 0.2000 2.0800 ;
        RECT 2.7600 1.6850 2.8500 2.0800 ;
        RECT 3.2800 1.6850 3.3700 2.0800 ;
        RECT 3.8000 1.6850 3.8900 2.0800 ;
        RECT 0.6400 1.6750 0.7300 2.0800 ;
        RECT 1.1650 1.6750 1.2550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.4100 0.9550 6.4650 1.0450 ;
      RECT 3.0200 0.4100 3.1100 0.8100 ;
      RECT 3.5400 0.4100 3.6300 0.8100 ;
      RECT 4.0600 0.4100 4.1500 0.8100 ;
      RECT 2.5600 0.8100 4.5000 0.9000 ;
      RECT 4.4100 0.9000 4.5000 0.9550 ;
      RECT 1.7150 1.4000 1.8050 1.7400 ;
      RECT 1.7150 1.3100 2.3300 1.4000 ;
      RECT 2.2400 1.4000 2.3300 1.7400 ;
      RECT 1.8550 0.9800 1.9450 1.3100 ;
      RECT 1.4650 0.8900 1.9450 0.9800 ;
      RECT 1.4650 0.5750 1.5550 0.8900 ;
      RECT 0.8500 0.4850 2.6500 0.5750 ;
      RECT 2.5600 0.5750 2.6500 0.8100 ;
      RECT 0.0550 1.2800 1.5600 1.3700 ;
      RECT 1.4700 1.2100 1.5600 1.2800 ;
      RECT 1.4700 1.1200 1.6800 1.2100 ;
      RECT 0.0550 0.9000 0.1450 1.2800 ;
      RECT 0.3700 1.3700 0.4600 1.8600 ;
      RECT 0.0550 0.8100 0.4600 0.9000 ;
      RECT 0.3700 0.4200 0.4600 0.8100 ;
      RECT 1.0100 0.9100 1.1000 1.2800 ;
      RECT 2.5000 1.2550 6.4650 1.2900 ;
      RECT 4.4350 1.2000 6.4650 1.2550 ;
      RECT 3.0200 1.3450 3.1100 1.7800 ;
      RECT 3.5400 1.3450 3.6300 1.7800 ;
      RECT 4.0600 1.3450 4.1500 1.7800 ;
      RECT 2.5000 1.2900 4.5250 1.3450 ;
      RECT 1.4250 1.8300 2.5900 1.9200 ;
      RECT 1.4250 1.5500 1.5150 1.8300 ;
      RECT 1.9750 1.4900 2.0650 1.8300 ;
      RECT 2.5000 1.3450 2.5900 1.8300 ;
      RECT 0.9050 1.4600 1.5150 1.5500 ;
      RECT 2.5000 1.1450 2.5900 1.2550 ;
      RECT 2.2850 1.0550 2.5900 1.1450 ;
      RECT 2.2850 0.7800 2.3750 1.0550 ;
      RECT 1.6450 0.6900 2.3750 0.7800 ;
      RECT 0.9050 1.5500 0.9950 1.8850 ;
  END
END BUFZ_X11M_A12TH

MACRO BUFZ_X16M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 10.0450 0.3200 ;
        RECT 0.1100 0.3200 0.2000 0.6300 ;
        RECT 0.6300 0.3200 0.7200 0.6100 ;
        RECT 1.1650 0.3200 1.2550 0.3900 ;
        RECT 3.2350 0.3200 3.4050 0.3950 ;
        RECT 3.7950 0.3200 3.8850 0.6450 ;
        RECT 4.3150 0.3200 4.4050 0.6550 ;
        RECT 4.8350 0.3200 4.9250 0.6550 ;
        RECT 5.3850 0.3200 5.4750 0.6300 ;
        RECT 5.8650 0.3200 6.0350 0.5250 ;
        RECT 6.3850 0.3200 6.5550 0.5250 ;
        RECT 6.9050 0.3200 7.0750 0.5250 ;
        RECT 7.4250 0.3200 7.5950 0.5250 ;
        RECT 7.9450 0.3200 8.1150 0.5250 ;
        RECT 8.4650 0.3200 8.6350 0.5250 ;
        RECT 8.9850 0.3200 9.1550 0.5250 ;
        RECT 9.5050 0.3200 9.6750 0.5250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 10.0450 2.7200 ;
        RECT 0.1100 1.7700 0.2000 2.0800 ;
        RECT 5.3850 1.7700 5.4750 2.0800 ;
        RECT 5.9050 1.7700 5.9950 2.0800 ;
        RECT 6.4250 1.7700 6.5150 2.0800 ;
        RECT 6.9450 1.7700 7.0350 2.0800 ;
        RECT 7.4650 1.7700 7.5550 2.0800 ;
        RECT 7.9850 1.7700 8.0750 2.0800 ;
        RECT 8.5050 1.7700 8.5950 2.0800 ;
        RECT 9.0250 1.7700 9.1150 2.0800 ;
        RECT 9.5450 1.7700 9.6350 2.0800 ;
        RECT 3.2750 1.6850 3.3650 2.0800 ;
        RECT 3.7950 1.6850 3.8850 2.0800 ;
        RECT 4.3150 1.6850 4.4050 2.0800 ;
        RECT 4.8350 1.6850 4.9250 2.0800 ;
        RECT 1.1250 1.6650 1.2950 2.0800 ;
        RECT 1.6450 1.6550 1.8150 2.0800 ;
        RECT 0.6400 1.5800 0.7300 2.0800 ;
    END
  END VDD

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3400 1.0500 0.7500 1.1500 ;
        RECT 0.6500 0.8000 0.7500 1.0500 ;
        RECT 0.6500 0.7000 1.8250 0.8000 ;
        RECT 1.7350 0.8000 1.8250 1.0200 ;
    END
    ANTENNAGATEAREA 0.51 ;
  END OE

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4950 1.0500 4.7150 1.1500 ;
    END
    ANTENNAGATEAREA 0.684 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6450 1.3900 9.8950 1.6100 ;
        RECT 5.6450 1.6100 5.7350 1.8200 ;
        RECT 6.1650 1.6100 6.2550 1.8200 ;
        RECT 6.6850 1.6100 6.7750 1.8200 ;
        RECT 7.2050 1.6100 7.2950 1.8200 ;
        RECT 7.7250 1.6100 7.8150 1.8200 ;
        RECT 8.2450 1.6100 8.3350 1.8200 ;
        RECT 8.7650 1.6100 8.8550 1.8200 ;
        RECT 9.2850 1.6100 9.3750 1.8200 ;
        RECT 9.8050 1.6100 9.8950 1.8200 ;
        RECT 9.3900 0.8400 9.6100 1.3900 ;
        RECT 5.6450 0.6200 9.8950 0.8400 ;
        RECT 5.6450 0.4250 5.7350 0.6200 ;
        RECT 6.1650 0.4250 6.2550 0.6200 ;
        RECT 6.6850 0.4250 6.7750 0.6200 ;
        RECT 7.2050 0.4250 7.2950 0.6200 ;
        RECT 7.7250 0.4250 7.8150 0.6200 ;
        RECT 8.2450 0.4250 8.3350 0.6200 ;
        RECT 8.7650 0.4250 8.8550 0.6200 ;
        RECT 9.2850 0.4250 9.3750 0.6200 ;
        RECT 9.8050 0.4250 9.8950 0.6200 ;
    END
    ANTENNADIFFAREA 2.6625 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0550 1.2550 1.9900 1.3450 ;
      RECT 1.9000 1.2100 1.9900 1.2550 ;
      RECT 1.9000 1.1200 2.1100 1.2100 ;
      RECT 1.1300 1.0000 1.2200 1.2550 ;
      RECT 0.9900 0.9100 1.2200 1.0000 ;
      RECT 0.0550 0.9000 0.1450 1.2550 ;
      RECT 0.3700 1.3450 0.4600 1.7200 ;
      RECT 0.0550 0.8100 0.4600 0.9000 ;
      RECT 0.3700 0.4900 0.4600 0.8100 ;
      RECT 3.0150 1.2550 8.8850 1.2700 ;
      RECT 5.3000 1.1800 8.8850 1.2550 ;
      RECT 0.9050 1.5450 0.9950 1.8850 ;
      RECT 1.4250 1.5450 1.5150 1.8850 ;
      RECT 1.9700 1.8300 3.1050 1.9200 ;
      RECT 1.9700 1.5450 2.0600 1.8300 ;
      RECT 2.4950 1.4900 2.5850 1.8300 ;
      RECT 3.0150 1.3450 3.1050 1.8300 ;
      RECT 0.9050 1.4550 2.0600 1.5450 ;
      RECT 3.0150 0.7800 3.1050 1.2550 ;
      RECT 2.1600 0.6900 3.1050 0.7800 ;
      RECT 3.5350 1.3450 3.6250 1.7800 ;
      RECT 4.0550 1.3450 4.1450 1.7800 ;
      RECT 4.5750 1.3450 4.6650 1.7800 ;
      RECT 5.0950 1.3450 5.1850 1.7800 ;
      RECT 3.0150 1.2700 5.3900 1.3450 ;
      RECT 5.2850 0.9500 8.8900 1.0400 ;
      RECT 2.2350 1.4000 2.3250 1.7400 ;
      RECT 2.2350 1.3100 2.8450 1.4000 ;
      RECT 2.7550 1.4000 2.8450 1.7400 ;
      RECT 2.2350 0.9800 2.3250 1.3100 ;
      RECT 1.9500 0.8900 2.3250 0.9800 ;
      RECT 1.9500 0.5750 2.0400 0.8900 ;
      RECT 0.8450 0.4850 3.6250 0.5750 ;
      RECT 3.5350 0.5750 3.6250 0.8100 ;
      RECT 4.0550 0.4100 4.1450 0.8100 ;
      RECT 4.5750 0.4100 4.6650 0.8100 ;
      RECT 3.5350 0.8100 5.3750 0.9000 ;
      RECT 5.2850 0.9000 5.3750 0.9500 ;
      RECT 5.0950 0.4100 5.1850 0.8100 ;
  END
END BUFZ_X16M_A12TH

MACRO BUFZ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.4300 0.3200 0.6000 0.7200 ;
        RECT 1.7100 0.3200 1.8000 0.6300 ;
    END
  END VSS

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0050 0.5550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END OE

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.6900 2.1500 1.4500 ;
        RECT 1.7900 1.4500 2.1500 1.5500 ;
        RECT 1.9100 0.6000 2.1500 0.6900 ;
        RECT 1.7900 1.5500 1.8800 1.8800 ;
    END
    ANTENNADIFFAREA 0.333125 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3400 1.0450 1.7250 1.1550 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.4300 1.4800 0.6000 2.0800 ;
        RECT 1.5300 1.4800 1.6200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0700 1.8800 0.3000 1.9700 ;
      RECT 0.2100 0.5000 0.3000 1.8800 ;
      RECT 0.0650 0.4100 0.3000 0.5000 ;
      RECT 0.7400 1.6650 1.3600 1.7550 ;
      RECT 1.2700 1.3700 1.3600 1.6650 ;
      RECT 1.1300 1.2800 1.3600 1.3700 ;
      RECT 1.0800 1.7550 1.1700 1.9650 ;
      RECT 0.7400 1.4600 0.8300 1.6650 ;
      RECT 1.1300 0.7800 1.2200 1.2800 ;
      RECT 0.9400 0.6900 1.2200 0.7800 ;
      RECT 1.3200 0.8000 1.9550 0.8900 ;
      RECT 1.8650 0.8900 1.9550 1.1600 ;
      RECT 0.7300 0.4800 1.4100 0.5700 ;
      RECT 1.3200 0.5700 1.4100 0.8000 ;
      RECT 0.9500 1.4850 1.1550 1.5750 ;
      RECT 0.9500 1.0500 1.0400 1.4850 ;
      RECT 0.7300 0.9600 1.0400 1.0500 ;
      RECT 0.7300 0.5700 0.8200 0.9600 ;
  END
END BUFZ_X1M_A12TH

MACRO BUFZ_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.5950 0.3200 0.6950 0.6300 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.0100 0.7500 1.1100 ;
        RECT 0.6450 1.1100 0.7500 1.2550 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END A

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.1850 1.9500 1.5050 ;
        RECT 1.2750 1.0500 1.9500 1.1850 ;
        RECT 1.2750 1.0150 1.3750 1.0500 ;
    END
    ANTENNAGATEAREA 0.0711 ;
  END OE

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.6200 0.4300 1.7500 ;
        RECT 0.3400 1.7500 0.4300 1.9900 ;
        RECT 0.0500 0.5850 0.1500 1.6200 ;
        RECT 0.0500 0.4950 0.4900 0.5850 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.0800 1.8400 0.1700 2.0800 ;
        RECT 1.7250 1.6050 1.8150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8550 0.5900 1.4600 0.6800 ;
      RECT 1.3700 0.6800 1.4600 0.8650 ;
      RECT 0.8550 1.6150 1.2400 1.7050 ;
      RECT 0.8550 0.9000 0.9500 1.6150 ;
      RECT 0.2750 0.8100 0.9500 0.9000 ;
      RECT 0.8550 0.6800 0.9500 0.8100 ;
      RECT 0.6500 1.8300 1.4750 1.9200 ;
      RECT 1.3850 1.4950 1.4750 1.8300 ;
      RECT 1.0950 1.4050 1.4750 1.4950 ;
      RECT 0.6500 1.4550 0.7400 1.8300 ;
      RECT 0.2650 1.3650 0.7400 1.4550 ;
      RECT 1.0950 0.7900 1.1850 1.4050 ;
      RECT 2.0250 1.7000 2.1500 1.9100 ;
      RECT 2.0600 0.7600 2.1500 1.7000 ;
      RECT 2.0250 0.6150 2.1500 0.7600 ;
      RECT 1.6350 0.5250 2.1500 0.6150 ;
      RECT 1.6350 0.5000 1.7500 0.5250 ;
      RECT 1.4300 0.4100 1.7500 0.5000 ;
  END
END BUFZ_X1P4M_A12TH

MACRO BUFZ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.7750 ;
        RECT 1.3400 0.3200 1.4300 0.3950 ;
        RECT 1.8750 0.3200 1.9650 0.3950 ;
        RECT 2.3950 0.3200 2.4850 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 2.0750 1.7700 2.1650 2.0800 ;
        RECT 2.6250 1.7700 2.7150 2.0800 ;
        RECT 0.4700 1.5300 0.5600 2.0800 ;
        RECT 1.3700 1.4400 1.4600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.9100 2.7500 1.4500 ;
        RECT 2.3650 1.4500 2.7500 1.5500 ;
        RECT 2.1350 0.8100 2.7500 0.9100 ;
        RECT 2.3650 1.5500 2.4550 1.8800 ;
        RECT 2.1350 0.4750 2.2250 0.8100 ;
    END
    ANTENNADIFFAREA 0.318 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3850 1.0500 1.8150 1.1500 ;
    END
    ANTENNAGATEAREA 0.105 ;
  END A

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8950 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0885 ;
  END OE
  OBS
    LAYER M1 ;
      RECT 0.0650 1.8800 0.3000 1.9700 ;
      RECT 0.2100 0.5100 0.3000 1.8800 ;
      RECT 0.0650 0.4200 0.3000 0.5100 ;
      RECT 1.9350 1.0300 2.1800 1.1200 ;
      RECT 1.9350 0.6050 2.0250 1.0300 ;
      RECT 0.7750 0.5150 2.0250 0.6050 ;
      RECT 1.5600 0.4100 1.7300 0.5150 ;
      RECT 0.7750 0.6050 0.8650 0.8950 ;
      RECT 0.7750 0.8950 1.0950 0.9850 ;
      RECT 1.0050 0.9850 1.0950 1.7200 ;
      RECT 1.1850 1.2400 2.5600 1.3300 ;
      RECT 2.4700 1.0400 2.5600 1.2400 ;
      RECT 0.7400 1.8300 1.2750 1.9200 ;
      RECT 0.7400 1.3800 0.8300 1.8300 ;
      RECT 1.1850 1.3300 1.2750 1.8300 ;
      RECT 1.1850 0.7850 1.2750 1.2400 ;
      RECT 0.9850 0.6950 1.2750 0.7850 ;
      RECT 1.6300 1.3300 1.7200 1.7400 ;
  END
END BUFZ_X2M_A12TH

MACRO BUFZ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.4700 0.3200 0.5600 0.6550 ;
        RECT 1.4150 0.3200 1.5050 0.4100 ;
        RECT 1.9750 0.3200 2.0650 0.4100 ;
        RECT 2.4950 0.3200 2.5850 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.0950 1.7700 2.1850 2.0800 ;
        RECT 2.6450 1.7700 2.7350 2.0800 ;
        RECT 1.4150 1.5800 1.5050 2.0800 ;
        RECT 0.4650 1.4850 0.5650 2.0800 ;
    END
  END VDD

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8600 0.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.1179 ;
  END OE

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4250 1.0450 1.8200 1.1550 ;
    END
    ANTENNAGATEAREA 0.144 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9500 3.1500 1.4500 ;
        RECT 2.3850 1.4500 3.1500 1.5500 ;
        RECT 2.2350 0.8500 3.1500 0.9500 ;
        RECT 2.3850 1.5500 2.4750 1.8800 ;
        RECT 2.9350 1.5500 3.0250 1.8800 ;
        RECT 2.2350 0.4700 2.3250 0.8500 ;
        RECT 2.7550 0.4700 2.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.64395 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2100 1.4450 0.3000 1.7650 ;
      RECT 0.0700 1.3550 0.3000 1.4450 ;
      RECT 0.0700 0.8350 0.1600 1.3550 ;
      RECT 0.0700 0.7450 0.3000 0.8350 ;
      RECT 0.2100 0.4400 0.3000 0.7450 ;
      RECT 0.6800 0.5150 2.1300 0.6050 ;
      RECT 2.0400 0.6050 2.1300 1.1500 ;
      RECT 1.0050 1.1750 1.0950 1.7400 ;
      RECT 0.6800 1.0850 1.0950 1.1750 ;
      RECT 0.6800 0.6050 0.7700 1.0850 ;
      RECT 1.2250 1.2600 2.9200 1.3500 ;
      RECT 2.8300 1.0400 2.9200 1.2600 ;
      RECT 0.7400 1.8300 1.3150 1.9200 ;
      RECT 0.7400 1.4900 0.8300 1.8300 ;
      RECT 1.2250 1.3500 1.3150 1.8300 ;
      RECT 1.2250 0.8150 1.3150 1.2600 ;
      RECT 0.9600 0.7250 1.3150 0.8150 ;
      RECT 1.6750 1.3500 1.7650 1.7400 ;
  END
END BUFZ_X3M_A12TH

MACRO BUFZ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.4300 0.3200 0.6000 0.6850 ;
        RECT 1.5200 0.3200 1.6100 0.4100 ;
        RECT 2.0800 0.3200 2.1700 0.4100 ;
        RECT 2.6000 0.3200 2.6900 0.6300 ;
        RECT 3.1200 0.3200 3.2100 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 1.5200 1.7700 1.6100 2.0800 ;
        RECT 2.1550 1.7700 2.2450 2.0800 ;
        RECT 2.7500 1.7700 2.8400 2.0800 ;
        RECT 3.2700 1.7700 3.3600 2.0800 ;
        RECT 0.4800 1.4900 0.5700 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.9500 3.5500 1.4500 ;
        RECT 2.4900 1.4500 3.5500 1.5500 ;
        RECT 2.3400 0.8500 3.5500 0.9500 ;
        RECT 2.4900 1.5500 2.5800 1.8800 ;
        RECT 3.0100 1.5500 3.1000 1.8800 ;
        RECT 2.3400 0.4700 2.4300 0.8500 ;
        RECT 2.8600 0.4700 2.9500 0.8500 ;
    END
    ANTENNADIFFAREA 0.636 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8950 1.8000 1.3050 ;
    END
    ANTENNAGATEAREA 0.1848 ;
  END A

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7750 0.5500 1.1950 ;
    END
    ANTENNAGATEAREA 0.1491 ;
  END OE
  OBS
    LAYER M1 ;
      RECT 0.2100 1.2900 0.9700 1.3800 ;
      RECT 0.8800 1.2100 0.9700 1.2900 ;
      RECT 0.8800 1.1200 1.2700 1.2100 ;
      RECT 0.2100 1.3800 0.3000 1.7300 ;
      RECT 0.2100 1.1000 0.3000 1.2900 ;
      RECT 0.0450 1.0100 0.3000 1.1000 ;
      RECT 0.2100 0.4100 0.3000 1.0100 ;
      RECT 0.7750 0.5000 2.2400 0.5900 ;
      RECT 2.1500 0.5900 2.2400 1.1450 ;
      RECT 1.0800 1.4200 1.1700 1.7400 ;
      RECT 1.0800 1.3300 1.4500 1.4200 ;
      RECT 1.3600 0.9500 1.4500 1.3300 ;
      RECT 0.7750 0.8600 1.4500 0.9500 ;
      RECT 0.7750 0.5900 0.8650 0.8600 ;
      RECT 1.9500 1.2600 3.2850 1.3500 ;
      RECT 3.1950 1.0400 3.2850 1.2600 ;
      RECT 1.3150 1.5500 2.0550 1.6400 ;
      RECT 1.7800 1.6400 1.8700 1.9600 ;
      RECT 1.9500 1.3500 2.0550 1.5500 ;
      RECT 1.9500 0.7700 2.0400 1.2600 ;
      RECT 0.9750 0.6800 2.0400 0.7700 ;
      RECT 0.8150 1.8300 1.4050 1.9200 ;
      RECT 1.3150 1.6400 1.4050 1.8300 ;
      RECT 0.8150 1.4900 0.9050 1.8300 ;
  END
END BUFZ_X4M_A12TH

MACRO BUFZ_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.4300 0.3200 0.6000 0.7000 ;
        RECT 2.0750 0.3200 2.1650 0.3950 ;
        RECT 2.5950 0.3200 2.6850 0.6100 ;
        RECT 3.0900 0.3200 3.2600 0.5050 ;
        RECT 3.6100 0.3200 3.7800 0.5050 ;
        RECT 4.1300 0.3200 4.3000 0.5050 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 2.0750 1.7700 2.1650 2.0800 ;
        RECT 2.6550 1.7700 2.7450 2.0800 ;
        RECT 3.2050 1.7700 3.2950 2.0800 ;
        RECT 3.7250 1.7700 3.8150 2.0800 ;
        RECT 4.2450 1.7700 4.3350 2.0800 ;
        RECT 0.4800 1.7100 0.5700 2.0800 ;
        RECT 1.0050 1.7100 1.0950 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0600 1.0500 2.5050 1.1500 ;
    END
    ANTENNAGATEAREA 0.2682 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.8200 4.5500 1.4500 ;
        RECT 2.9450 1.4500 4.5950 1.5500 ;
        RECT 2.8700 0.7200 4.5500 0.8200 ;
        RECT 2.9450 1.5500 3.0350 1.8800 ;
        RECT 3.4650 1.5500 3.5550 1.8800 ;
        RECT 3.9850 1.5500 4.0750 1.8800 ;
        RECT 4.5050 1.5500 4.5950 1.8800 ;
        RECT 2.8700 0.4100 2.9600 0.7200 ;
        RECT 3.3900 0.4100 3.4800 0.7200 ;
        RECT 3.9100 0.4100 4.0000 0.7200 ;
        RECT 4.4600 0.4100 4.5500 0.7200 ;
    END
    ANTENNADIFFAREA 1.054 ;
  END Y

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9500 0.5500 1.2500 ;
        RECT 0.4500 0.8500 1.1900 0.9500 ;
        RECT 1.1000 0.9500 1.1900 1.1350 ;
    END
    ANTENNAGATEAREA 0.2082 ;
  END OE
  OBS
    LAYER M1 ;
      RECT 0.2100 1.3400 1.2850 1.4300 ;
      RECT 1.1950 1.2250 1.2850 1.3400 ;
      RECT 0.8300 1.0800 0.9200 1.3400 ;
      RECT 0.2100 1.4300 0.3000 1.7600 ;
      RECT 0.2100 0.5400 0.3000 1.3400 ;
      RECT 1.8150 1.2600 4.1200 1.3500 ;
      RECT 0.7450 1.6100 0.8350 1.9900 ;
      RECT 1.2900 1.8300 1.9050 1.9200 ;
      RECT 1.2900 1.6100 1.3800 1.8300 ;
      RECT 1.8150 1.3500 1.9050 1.8300 ;
      RECT 0.7450 1.5200 1.3800 1.6100 ;
      RECT 1.8150 0.7800 1.9050 1.2600 ;
      RECT 1.4800 0.6900 1.9050 0.7800 ;
      RECT 2.3350 1.3500 2.4250 1.7400 ;
      RECT 2.6850 0.9300 4.1200 1.0200 ;
      RECT 0.6900 0.4850 2.5050 0.5750 ;
      RECT 2.4150 0.5750 2.5050 0.7200 ;
      RECT 1.5550 0.9600 1.6450 1.7100 ;
      RECT 1.2800 0.8700 1.6450 0.9600 ;
      RECT 1.2800 0.5750 1.3700 0.8700 ;
      RECT 2.4150 0.7200 2.7750 0.8100 ;
      RECT 2.6850 0.8100 2.7750 0.9300 ;
  END
END BUFZ_X6M_A12TH

MACRO BUFZ_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.6600 ;
        RECT 1.9600 0.3200 2.0500 0.3950 ;
        RECT 2.4800 0.3200 2.5700 0.6300 ;
        RECT 3.0300 0.3200 3.1200 0.6300 ;
        RECT 3.5100 0.3200 3.6800 0.5200 ;
        RECT 4.0300 0.3200 4.2000 0.5200 ;
        RECT 4.5500 0.3200 4.7200 0.5200 ;
        RECT 5.0700 0.3200 5.2400 0.5200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.3700 1.7700 0.4600 2.0800 ;
        RECT 0.8900 1.7700 0.9800 2.0800 ;
        RECT 1.9600 1.7700 2.0500 2.0800 ;
        RECT 2.4800 1.7700 2.5700 2.0800 ;
        RECT 3.0600 1.7700 3.1500 2.0800 ;
        RECT 3.5800 1.7700 3.6700 2.0800 ;
        RECT 4.1000 1.7700 4.1900 2.0800 ;
        RECT 4.6200 1.7700 4.7100 2.0800 ;
        RECT 5.1400 1.7700 5.2300 2.0800 ;
    END
  END VDD

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.1000 0.5550 1.1900 ;
        RECT 0.4450 0.9500 0.5550 1.1000 ;
        RECT 0.4450 0.8500 1.1050 0.9500 ;
    END
    ANTENNAGATEAREA 0.2574 ;
  END OE

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8800 1.0500 2.6150 1.1500 ;
    END
    ANTENNAGATEAREA 0.348 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3200 1.4350 5.4900 1.5650 ;
        RECT 3.3200 1.5650 3.4100 1.8700 ;
        RECT 3.8400 1.5650 3.9300 1.8700 ;
        RECT 4.3600 1.5650 4.4500 1.8700 ;
        RECT 4.8800 1.5650 4.9700 1.8700 ;
        RECT 5.4000 1.5650 5.4900 1.8700 ;
        RECT 5.2350 0.8300 5.3650 1.4350 ;
        RECT 3.2900 0.7000 5.4600 0.8300 ;
        RECT 3.2900 0.4200 3.3800 0.7000 ;
        RECT 3.8100 0.4200 3.9000 0.7000 ;
        RECT 4.3300 0.4200 4.4200 0.7000 ;
        RECT 4.8500 0.4200 4.9400 0.7000 ;
        RECT 5.3700 0.4200 5.4600 0.7000 ;
    END
    ANTENNADIFFAREA 1.3845 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0950 1.2800 1.2850 1.3700 ;
      RECT 1.1950 1.0900 1.2850 1.2800 ;
      RECT 0.7350 1.0400 0.8250 1.2800 ;
      RECT 0.0950 1.3700 0.1850 1.7200 ;
      RECT 0.0950 0.5000 0.1850 1.2800 ;
      RECT 3.1000 1.2100 4.8700 1.3000 ;
      RECT 0.6300 1.5500 0.7200 1.8700 ;
      RECT 1.1750 1.8300 1.7900 1.9200 ;
      RECT 1.1750 1.5500 1.2650 1.8300 ;
      RECT 1.7000 1.4400 1.7900 1.8300 ;
      RECT 0.6300 1.4600 1.2650 1.5500 ;
      RECT 1.7000 0.7800 1.7900 1.3500 ;
      RECT 1.3750 0.6900 1.7900 0.7800 ;
      RECT 2.2200 1.4400 2.3100 1.7800 ;
      RECT 2.7400 1.4400 2.8300 1.7800 ;
      RECT 1.7000 1.3500 3.1900 1.4400 ;
      RECT 3.1000 1.3000 3.1900 1.3500 ;
      RECT 3.1100 0.9400 4.9000 1.0300 ;
      RECT 0.5700 0.4850 2.3900 0.5750 ;
      RECT 2.3000 0.5750 2.3900 0.8100 ;
      RECT 1.4400 1.0000 1.5300 1.7400 ;
      RECT 1.1950 0.9100 1.5300 1.0000 ;
      RECT 1.1950 0.5750 1.2850 0.9100 ;
      RECT 2.7400 0.4200 2.8300 0.8100 ;
      RECT 2.3000 0.8100 3.2000 0.9000 ;
      RECT 3.1100 0.9000 3.2000 0.9400 ;
  END
END BUFZ_X8M_A12TH

MACRO AOI31_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1000 0.3200 0.1900 0.6300 ;
        RECT 1.6200 0.3200 1.7900 0.5200 ;
        RECT 3.1800 0.3200 3.3500 0.5200 ;
        RECT 3.8150 0.3200 3.9050 0.7600 ;
        RECT 4.3350 0.3200 4.4250 0.7950 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 1.2500 2.0850 1.3500 ;
        RECT 1.3150 1.2100 1.4050 1.2500 ;
        RECT 1.9950 1.2100 2.0850 1.2500 ;
        RECT 1.2050 1.0600 1.4050 1.2100 ;
        RECT 1.9950 1.0600 2.2050 1.2100 ;
        RECT 0.5150 0.9700 1.4050 1.0600 ;
        RECT 1.9950 0.9700 2.9450 1.0600 ;
        RECT 0.5150 1.0600 0.6050 1.2400 ;
        RECT 2.8550 1.0600 2.9450 1.2400 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8800 1.7500 1.0700 ;
        RECT 1.5150 1.0700 1.8850 1.1600 ;
        RECT 0.2550 0.7900 3.2050 0.8800 ;
        RECT 0.2550 0.8800 0.3450 1.2400 ;
        RECT 3.1150 0.8800 3.2050 1.2400 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6100 1.0500 4.0900 1.1500 ;
    END
    ANTENNAGATEAREA 0.2916 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.2500 1.1050 1.3500 ;
        RECT 1.0150 1.3500 1.1050 1.4400 ;
        RECT 0.7350 1.1500 1.1050 1.2500 ;
        RECT 1.0150 1.4400 2.3850 1.5300 ;
        RECT 2.2950 1.2400 2.3850 1.4400 ;
        RECT 2.2950 1.1500 2.7150 1.2400 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4000 0.8500 4.1700 0.9500 ;
        RECT 3.4000 0.9500 3.5000 1.3000 ;
        RECT 3.4000 0.7000 3.6450 0.8500 ;
        RECT 4.0700 0.4100 4.1700 0.8500 ;
        RECT 3.4000 1.3000 4.1700 1.3900 ;
        RECT 0.8400 0.6100 3.6450 0.7000 ;
        RECT 3.5500 1.3900 3.6500 1.7150 ;
        RECT 4.0700 1.3900 4.1700 1.7150 ;
        RECT 0.8400 0.4100 1.0100 0.6100 ;
        RECT 2.4000 0.4100 2.5700 0.6100 ;
        RECT 3.5550 0.4100 3.6450 0.6100 ;
    END
    ANTENNADIFFAREA 0.794 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.3600 1.8000 0.4500 2.0800 ;
        RECT 0.8800 1.8000 0.9700 2.0800 ;
        RECT 1.4000 1.8000 1.4900 2.0800 ;
        RECT 1.9200 1.8000 2.0100 2.0800 ;
        RECT 2.4400 1.8000 2.5300 2.0800 ;
        RECT 3.0050 1.8000 3.0950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.2950 1.8300 4.4250 1.9200 ;
      RECT 4.3350 1.5100 4.4250 1.8300 ;
      RECT 0.1000 1.6200 3.3850 1.7100 ;
      RECT 3.2950 1.7100 3.3850 1.8300 ;
      RECT 3.2950 1.5300 3.3850 1.6200 ;
      RECT 3.8150 1.5100 3.9050 1.8300 ;
      RECT 0.1000 1.7100 0.1900 1.9900 ;
      RECT 0.6200 1.7100 0.7100 1.9900 ;
      RECT 1.1400 1.7100 1.2300 1.9900 ;
      RECT 1.6600 1.7100 1.7500 1.9900 ;
      RECT 2.1800 1.7100 2.2700 1.9900 ;
      RECT 2.7000 1.7100 2.7900 1.9900 ;
  END
END AOI31_X4M_A12TH

MACRO AOI31_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6350 ;
        RECT 1.6000 0.3200 1.7700 0.5200 ;
        RECT 3.2100 0.3200 3.3800 0.5200 ;
        RECT 4.7700 0.3200 4.9400 0.5200 ;
        RECT 5.4050 0.3200 5.4950 0.6000 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3050 1.2500 2.0550 1.3500 ;
        RECT 1.9650 1.2100 2.0550 1.2500 ;
        RECT 1.3050 1.2100 1.3950 1.2500 ;
        RECT 1.9650 1.0600 2.1750 1.2100 ;
        RECT 1.1850 1.0600 1.3950 1.2100 ;
        RECT 1.9650 0.9700 3.0150 1.0600 ;
        RECT 0.4950 0.9700 1.3950 1.0600 ;
        RECT 2.8050 1.0600 3.0150 1.2100 ;
        RECT 0.4950 1.0600 0.5850 1.2400 ;
        RECT 2.9250 1.2100 3.0150 1.2600 ;
        RECT 2.9250 1.2600 3.6650 1.3500 ;
        RECT 3.5750 1.2100 3.6650 1.2600 ;
        RECT 3.5750 1.0600 3.7850 1.2100 ;
        RECT 3.5750 0.9700 4.5350 1.0600 ;
        RECT 4.4450 1.0600 4.5350 1.2400 ;
    END
    ANTENNAGATEAREA 0.5868 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8800 1.8750 1.0700 ;
        RECT 1.5050 1.0700 1.8750 1.1600 ;
        RECT 0.2350 0.7900 3.1950 0.8800 ;
        RECT 0.2350 0.8800 0.3250 1.2400 ;
        RECT 3.1050 0.8800 3.1950 1.0800 ;
        RECT 3.1050 1.0800 3.4850 1.1700 ;
        RECT 3.3950 0.8800 3.4850 1.0800 ;
        RECT 3.3950 0.7900 4.7950 0.8800 ;
        RECT 4.7050 0.8800 4.7950 1.2400 ;
    END
    ANTENNAGATEAREA 0.5868 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.2500 1.0850 1.3500 ;
        RECT 0.9950 1.3500 1.0850 1.4400 ;
        RECT 0.7150 1.1500 1.0850 1.2500 ;
        RECT 0.9950 1.4400 3.9650 1.5300 ;
        RECT 2.5850 1.2400 2.6750 1.4400 ;
        RECT 3.8750 1.2400 3.9650 1.4400 ;
        RECT 2.3050 1.1500 2.6750 1.2400 ;
        RECT 3.8750 1.1500 4.2850 1.2400 ;
    END
    ANTENNAGATEAREA 0.5868 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2050 1.0600 6.2050 1.1600 ;
        RECT 5.6100 1.0500 5.7900 1.0600 ;
    END
    ANTENNAGATEAREA 0.4374 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9950 1.2500 6.2650 1.3400 ;
        RECT 5.1250 1.3400 6.2650 1.3500 ;
        RECT 4.9950 0.7800 5.0950 1.2500 ;
        RECT 5.1250 1.3500 5.2250 1.7400 ;
        RECT 5.6450 1.3500 5.7450 1.7400 ;
        RECT 6.1650 1.3500 6.2650 1.7400 ;
        RECT 4.9950 0.7000 5.7600 0.7800 ;
        RECT 0.8200 0.6900 5.7600 0.7000 ;
        RECT 0.8200 0.6100 5.2400 0.6900 ;
        RECT 5.6600 0.4100 5.7600 0.6900 ;
        RECT 0.8200 0.4100 0.9900 0.6100 ;
        RECT 2.4000 0.4100 2.5700 0.6100 ;
        RECT 3.9900 0.4100 4.1600 0.6100 ;
        RECT 5.1400 0.4100 5.2400 0.6100 ;
    END
    ANTENNADIFFAREA 1.2863 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.3400 1.8000 0.4300 2.0800 ;
        RECT 0.8600 1.8000 0.9500 2.0800 ;
        RECT 1.3800 1.8000 1.4700 2.0800 ;
        RECT 1.9000 1.8000 1.9900 2.0800 ;
        RECT 2.4500 1.8000 2.5400 2.0800 ;
        RECT 2.9900 1.8000 3.0800 2.0800 ;
        RECT 3.5100 1.8000 3.6000 2.0800 ;
        RECT 4.0300 1.8000 4.1200 2.0800 ;
        RECT 4.5900 1.8000 4.6800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.8700 1.8300 6.5200 1.9200 ;
      RECT 6.4300 1.4900 6.5200 1.8300 ;
      RECT 0.0800 1.6200 4.9600 1.7100 ;
      RECT 4.8700 1.7100 4.9600 1.8300 ;
      RECT 4.8700 1.5500 4.9600 1.6200 ;
      RECT 5.3900 1.4900 5.4800 1.8300 ;
      RECT 5.9100 1.4900 6.0000 1.8300 ;
      RECT 0.0800 1.7100 0.1700 1.9900 ;
      RECT 0.6000 1.7100 0.6900 1.9900 ;
      RECT 1.1200 1.7100 1.2100 1.9900 ;
      RECT 1.6400 1.7100 1.7300 1.9900 ;
      RECT 2.1600 1.7100 2.2500 1.9900 ;
      RECT 2.7300 1.7100 2.8200 1.9900 ;
      RECT 3.2500 1.7100 3.3400 1.9900 ;
      RECT 3.7700 1.7100 3.8600 1.9900 ;
      RECT 4.2900 1.7100 4.3800 1.9900 ;
  END
END AOI31_X6M_A12TH

MACRO AOI32_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7200 ;
        RECT 1.4100 0.3200 1.5100 0.5200 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 0.8500 0.9150 0.9500 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.2500 0.7100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.7950 0.3600 1.1550 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9700 1.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0426 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7000 1.5500 1.6100 ;
        RECT 1.1150 1.6100 1.5500 1.7100 ;
        RECT 0.7800 0.6100 1.5500 0.7000 ;
        RECT 0.7800 0.4100 0.9500 0.6100 ;
    END
    ANTENNADIFFAREA 0.181375 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8100 1.3500 1.2300 ;
    END
    ANTENNAGATEAREA 0.0426 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.6200 1.6650 0.7200 2.0800 ;
        RECT 0.0900 1.6000 0.1900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8550 1.8200 1.5450 1.9200 ;
      RECT 0.8550 1.5750 1.0250 1.8200 ;
      RECT 0.3500 1.4850 1.0250 1.5750 ;
      RECT 0.3500 1.5750 0.4500 1.9900 ;
  END
END AOI32_X0P5M_A12TH

MACRO AOI32_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6500 ;
        RECT 1.4100 0.3200 1.5100 0.4550 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 0.8500 0.9100 0.9600 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.2500 0.7100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.7450 0.3550 1.1450 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.0400 1.1500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7000 1.5500 1.6100 ;
        RECT 1.0950 1.6100 1.5500 1.7100 ;
        RECT 0.7800 0.6100 1.5500 0.7000 ;
        RECT 0.7800 0.4100 0.9500 0.6100 ;
    END
    ANTENNADIFFAREA 0.256875 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8900 1.3500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0603 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.6200 1.6900 0.7200 2.0800 ;
        RECT 0.0900 1.6800 0.1900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8950 1.8300 1.5450 1.9200 ;
      RECT 0.8950 1.6000 0.9850 1.8300 ;
      RECT 0.3550 1.5100 0.9850 1.6000 ;
      RECT 0.3550 1.6000 0.4450 1.9500 ;
  END
END AOI32_X0P7M_A12TH

MACRO AOI32_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6250 ;
        RECT 1.3750 0.3200 1.5450 0.5200 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.1000 0.8700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8900 0.5500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.0800 0.3500 1.3200 ;
        RECT 0.2500 0.8900 0.3500 1.0800 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8150 1.1500 1.2350 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7000 1.5500 1.6100 ;
        RECT 1.0950 1.6100 1.5500 1.7100 ;
        RECT 0.8550 0.6100 1.5500 0.7000 ;
        RECT 0.8550 0.4100 1.0250 0.6100 ;
    END
    ANTENNADIFFAREA 0.31375 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9700 1.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6200 1.7700 0.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8800 1.8200 1.5450 1.9200 ;
      RECT 0.8800 1.5900 0.9800 1.8200 ;
      RECT 0.3500 1.5000 0.9800 1.5900 ;
      RECT 0.3500 1.5900 0.4500 1.9200 ;
  END
END AOI32_X1M_A12TH

MACRO AOI32_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.0850 0.3200 0.1950 0.7950 ;
        RECT 1.6850 0.3200 1.8550 0.7100 ;
        RECT 2.7450 0.3200 2.9150 0.7000 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.2450 1.1200 1.3550 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.3200 0.5500 1.6500 ;
        RECT 0.4500 1.6500 1.4050 1.7400 ;
        RECT 1.3050 1.3300 1.4050 1.6500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 1.6600 1.1000 ;
        RECT 0.2400 1.1000 0.3500 1.2300 ;
        RECT 1.5600 1.1000 1.6600 1.1800 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0950 1.2500 2.5050 1.3600 ;
    END
    ANTENNAGATEAREA 0.1206 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.9000 2.9500 1.6400 ;
        RECT 1.9250 1.6400 2.9500 1.7400 ;
        RECT 0.9050 0.8000 2.9500 0.9000 ;
        RECT 0.9050 0.7000 1.0050 0.8000 ;
        RECT 2.2550 0.5300 2.3650 0.8000 ;
    END
    ANTENNADIFFAREA 0.46055 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0500 2.7250 1.1500 ;
        RECT 2.6250 1.1500 2.7250 1.2400 ;
    END
    ANTENNAGATEAREA 0.1206 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.3650 2.0100 0.4750 2.0800 ;
        RECT 0.9000 2.0100 1.0100 2.0800 ;
        RECT 1.4550 2.0100 1.5650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.8300 2.9350 1.9200 ;
  END
END AOI32_X1P4M_A12TH

MACRO AOI32_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.1100 0.3200 0.2100 0.6300 ;
        RECT 1.6850 0.3200 1.8550 0.5500 ;
        RECT 2.7450 0.3200 2.9150 0.5500 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2400 0.3500 1.4900 ;
        RECT 0.2500 1.4900 1.6650 1.5800 ;
        RECT 0.2100 1.0700 0.3500 1.2400 ;
        RECT 1.5650 1.0700 1.6650 1.4900 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7600 0.5600 1.2350 ;
        RECT 0.4500 0.6700 1.3850 0.7600 ;
        RECT 1.2850 0.7600 1.3850 1.2400 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.0500 1.1100 1.2000 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0950 1.0500 2.5050 1.1600 ;
    END
    ANTENNAGATEAREA 0.1704 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6300 1.0800 2.7500 1.3900 ;
        RECT 1.8200 1.3900 2.7500 1.4900 ;
        RECT 1.8200 1.0700 1.9200 1.3900 ;
    END
    ANTENNAGATEAREA 0.1704 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.3700 2.0100 0.4700 2.0800 ;
        RECT 0.8900 2.0100 0.9900 2.0800 ;
        RECT 1.4600 2.0100 1.5600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.7600 2.9500 1.6200 ;
        RECT 1.9250 1.6200 2.9500 1.7200 ;
        RECT 1.4950 0.6600 2.9500 0.7600 ;
        RECT 1.4950 0.5700 1.5950 0.6600 ;
        RECT 2.2500 0.5250 2.3500 0.6600 ;
        RECT 0.8500 0.4800 1.5950 0.5700 ;
    END
    ANTENNADIFFAREA 0.6443 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0550 1.8200 2.9350 1.9200 ;
  END
END AOI32_X2M_A12TH

MACRO AOI32_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.6100 0.3200 0.7100 0.6300 ;
        RECT 3.4700 0.3200 3.5700 0.7700 ;
        RECT 4.0100 0.3200 4.1100 0.8400 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8800 1.0500 2.3200 1.1600 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0800 1.0500 1.5200 1.1600 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0500 0.7200 1.1600 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6800 1.0500 3.1200 1.1600 ;
    END
    ANTENNAGATEAREA 0.2556 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9550 2.5500 1.2800 ;
        RECT 2.4500 1.2800 3.8350 1.3800 ;
        RECT 1.9100 0.8650 3.0500 0.9550 ;
        RECT 2.6900 1.3800 2.7900 1.7400 ;
        RECT 3.2100 1.3800 3.3100 1.7400 ;
        RECT 3.7350 1.3800 3.8350 1.7400 ;
        RECT 1.9100 0.7450 2.0100 0.8650 ;
        RECT 2.9500 0.7450 3.0500 0.8650 ;
        RECT 2.4300 0.5250 2.5300 0.8650 ;
    END
    ANTENNADIFFAREA 0.93535 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4800 1.0500 3.9200 1.1600 ;
    END
    ANTENNAGATEAREA 0.2556 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 0.8700 1.4850 0.9600 ;
      RECT 1.3950 0.7500 1.4850 0.8700 ;
      RECT 0.8750 0.5300 0.9650 0.8700 ;
      RECT 0.3550 0.5300 0.4450 0.8700 ;
      RECT 1.0950 0.4800 2.3050 0.5700 ;
      RECT 2.1350 0.5700 2.3050 0.7700 ;
      RECT 1.0950 0.5700 1.2650 0.7800 ;
      RECT 1.6550 0.5700 1.7450 0.9100 ;
      RECT 3.2150 0.8600 3.8350 0.9500 ;
      RECT 3.7450 0.5200 3.8350 0.8600 ;
      RECT 3.2150 0.5700 3.3050 0.8600 ;
      RECT 2.6550 0.4800 3.3050 0.5700 ;
      RECT 2.6550 0.5700 2.8250 0.7700 ;
      RECT 2.4350 1.8300 4.1050 1.9200 ;
      RECT 4.0150 1.4900 4.1050 1.8300 ;
      RECT 0.3550 1.4900 2.5250 1.5800 ;
      RECT 2.4350 1.5800 2.5250 1.8300 ;
      RECT 2.9550 1.4900 3.0450 1.8300 ;
      RECT 3.4750 1.4900 3.5650 1.8300 ;
      RECT 0.3550 1.5800 0.4450 1.9200 ;
      RECT 0.8750 1.5800 0.9650 1.9200 ;
      RECT 1.3950 1.5800 1.4850 1.9200 ;
      RECT 1.9150 1.5800 2.0050 1.9200 ;
  END
END AOI32_X3M_A12TH

MACRO AOI32_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1800 0.6300 ;
        RECT 1.6100 0.3200 1.7800 0.5200 ;
        RECT 3.1700 0.3200 3.3400 0.5200 ;
        RECT 4.3400 0.3200 4.4300 0.5800 ;
        RECT 5.4300 0.3200 5.5200 0.6500 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 1.2500 2.0650 1.3500 ;
        RECT 1.3150 1.2100 1.4050 1.2500 ;
        RECT 1.9750 1.2100 2.0650 1.2500 ;
        RECT 1.1950 1.0600 1.4050 1.2100 ;
        RECT 1.9750 1.0600 2.1650 1.2100 ;
        RECT 0.5050 0.9700 1.4050 1.0600 ;
        RECT 1.9750 0.9700 2.9350 1.0600 ;
        RECT 0.5050 1.0600 0.5950 1.2400 ;
        RECT 2.8450 1.0600 2.9350 1.2400 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8800 1.8850 1.0700 ;
        RECT 1.5150 1.0700 1.8850 1.1600 ;
        RECT 0.2450 0.7900 3.1650 0.8800 ;
        RECT 0.2450 0.8800 0.3350 1.2400 ;
        RECT 3.0750 0.8800 3.1650 1.2600 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6100 0.8700 5.1350 0.9600 ;
        RECT 3.6100 0.8600 4.0450 0.8700 ;
        RECT 3.6100 0.8500 3.7900 0.8600 ;
    END
    ANTENNAGATEAREA 0.3408 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.2500 1.0950 1.3500 ;
        RECT 1.0050 1.3500 1.0950 1.4400 ;
        RECT 0.7250 1.1500 1.0950 1.2500 ;
        RECT 1.0050 1.4400 2.3450 1.5300 ;
        RECT 2.2550 1.2400 2.3450 1.4400 ;
        RECT 2.2550 1.1500 2.6350 1.2400 ;
    END
    ANTENNAGATEAREA 0.3912 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4350 1.0500 5.4700 1.1400 ;
        RECT 4.2000 1.1400 4.5700 1.1500 ;
    END
    ANTENNAGATEAREA 0.3408 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2550 1.2600 5.2150 1.3500 ;
        RECT 3.5550 1.3500 3.6550 1.7300 ;
        RECT 4.0750 1.3500 4.1750 1.7300 ;
        RECT 4.5950 1.3500 4.6950 1.7300 ;
        RECT 5.1150 1.3500 5.2150 1.7300 ;
        RECT 3.5600 1.2500 5.2150 1.2600 ;
        RECT 3.2550 0.7600 3.3450 1.2600 ;
        RECT 3.2550 0.7000 4.9900 0.7600 ;
        RECT 0.8300 0.6700 4.9900 0.7000 ;
        RECT 0.8300 0.6100 3.3450 0.6700 ;
        RECT 3.7800 0.4300 3.9500 0.6700 ;
        RECT 4.8200 0.4300 4.9900 0.6700 ;
        RECT 0.8300 0.4100 1.0000 0.6100 ;
        RECT 2.3900 0.4100 2.5600 0.6100 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.3500 1.8000 0.4400 2.0800 ;
        RECT 0.8700 1.8000 0.9600 2.0800 ;
        RECT 1.3900 1.8000 1.4800 2.0800 ;
        RECT 1.9100 1.8000 2.0000 2.0800 ;
        RECT 2.4300 1.8000 2.5200 2.0800 ;
        RECT 2.9950 1.8000 3.0850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.3000 1.8300 5.4700 1.9200 ;
      RECT 5.3800 1.4850 5.4700 1.8300 ;
      RECT 0.0900 1.6200 3.3900 1.7100 ;
      RECT 3.3000 1.7100 3.3900 1.8300 ;
      RECT 3.3000 1.5500 3.3900 1.6200 ;
      RECT 3.8200 1.4850 3.9100 1.8300 ;
      RECT 4.3400 1.4850 4.4300 1.8300 ;
      RECT 4.8600 1.4850 4.9500 1.8300 ;
      RECT 0.0900 1.7100 0.1800 1.9900 ;
      RECT 0.6100 1.7100 0.7000 1.9900 ;
      RECT 1.1300 1.7100 1.2200 1.9900 ;
      RECT 1.6500 1.7100 1.7400 1.9900 ;
      RECT 2.1700 1.7100 2.2600 1.9900 ;
      RECT 2.6900 1.7100 2.7800 1.9900 ;
  END
END AOI32_X4M_A12TH

MACRO AOI32_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6300 ;
        RECT 1.6000 0.3200 1.7700 0.5200 ;
        RECT 3.1600 0.3200 3.3300 0.5200 ;
        RECT 4.7200 0.3200 4.8900 0.5200 ;
        RECT 5.9300 0.3200 6.0200 0.5800 ;
        RECT 6.9700 0.3200 7.0600 0.5800 ;
        RECT 8.0100 0.3200 8.1000 0.6500 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3050 1.2500 2.0750 1.3500 ;
        RECT 1.9850 1.2100 2.0750 1.2500 ;
        RECT 1.3050 1.2100 1.3950 1.2500 ;
        RECT 1.9850 1.0600 2.1750 1.2100 ;
        RECT 1.1850 1.0600 1.3950 1.2100 ;
        RECT 1.9850 0.9700 2.9650 1.0600 ;
        RECT 0.4950 0.9700 1.3950 1.0600 ;
        RECT 2.7550 1.0600 2.9650 1.2100 ;
        RECT 0.4950 1.0600 0.5850 1.2400 ;
        RECT 2.8750 1.2100 2.9650 1.2600 ;
        RECT 2.8750 1.2600 3.6050 1.3500 ;
        RECT 3.5150 1.2100 3.6050 1.2600 ;
        RECT 3.5150 1.0600 3.7150 1.2100 ;
        RECT 3.5150 0.9700 4.4850 1.0600 ;
        RECT 4.3950 1.0600 4.4850 1.2400 ;
    END
    ANTENNAGATEAREA 0.5868 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8800 1.7500 1.0700 ;
        RECT 0.3150 0.7900 3.1450 0.8800 ;
        RECT 1.5050 1.0700 1.8750 1.1600 ;
        RECT 0.3150 0.8800 0.4050 1.0300 ;
        RECT 3.0550 0.8800 3.1450 1.0800 ;
        RECT 0.2350 1.0300 0.4050 1.1200 ;
        RECT 3.0550 1.0800 3.4250 1.1700 ;
        RECT 0.2350 1.1200 0.3250 1.2400 ;
        RECT 3.3350 0.8800 3.4250 1.0800 ;
        RECT 3.3350 0.7900 4.7150 0.8800 ;
        RECT 4.6250 0.8800 4.7150 1.2600 ;
    END
    ANTENNAGATEAREA 0.5868 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3200 0.8900 7.7150 0.9600 ;
        RECT 5.3200 0.9600 5.6300 0.9800 ;
        RECT 6.3050 0.9600 7.7150 0.9800 ;
        RECT 5.3200 0.8700 6.3950 0.8900 ;
        RECT 5.3200 0.8500 5.5900 0.8700 ;
    END
    ANTENNAGATEAREA 0.5112 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.2500 1.0850 1.3500 ;
        RECT 0.9950 1.3500 1.0850 1.4400 ;
        RECT 0.7150 1.1500 1.0850 1.2500 ;
        RECT 0.9950 1.4400 3.8950 1.5300 ;
        RECT 2.5550 1.2400 2.6450 1.4400 ;
        RECT 3.8050 1.2400 3.8950 1.4400 ;
        RECT 2.2850 1.1500 2.6450 1.2400 ;
        RECT 3.8050 1.1500 4.2050 1.2400 ;
    END
    ANTENNAGATEAREA 0.5868 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0050 1.0700 8.0250 1.1600 ;
        RECT 5.7200 1.0600 6.1550 1.0700 ;
        RECT 5.8100 1.0500 5.9900 1.0600 ;
    END
    ANTENNAGATEAREA 0.5112 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8050 1.2500 7.8400 1.3400 ;
        RECT 5.1500 1.3400 7.8400 1.3500 ;
        RECT 4.8050 0.7600 4.8950 1.2500 ;
        RECT 5.1500 1.3500 5.2400 1.7400 ;
        RECT 5.6700 1.3500 5.7600 1.7400 ;
        RECT 6.1900 1.3500 6.2800 1.7400 ;
        RECT 6.7100 1.3500 6.8000 1.7400 ;
        RECT 7.2300 1.3500 7.3200 1.7400 ;
        RECT 7.7500 1.3500 7.8400 1.7400 ;
        RECT 4.8050 0.7000 7.5800 0.7600 ;
        RECT 6.4500 0.7600 6.5400 0.7800 ;
        RECT 7.4900 0.7600 7.5800 0.7800 ;
        RECT 0.8200 0.6700 7.5800 0.7000 ;
        RECT 0.8200 0.6100 4.8950 0.6700 ;
        RECT 5.3700 0.4500 5.5400 0.6700 ;
        RECT 6.4500 0.4100 6.5400 0.6700 ;
        RECT 7.4900 0.4100 7.5800 0.6700 ;
        RECT 0.8200 0.4100 0.9900 0.6100 ;
        RECT 2.3800 0.4100 2.5500 0.6100 ;
        RECT 3.9400 0.4100 4.1100 0.6100 ;
    END
    ANTENNADIFFAREA 1.83 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 0.3400 1.8000 0.4300 2.0800 ;
        RECT 0.8600 1.8000 0.9500 2.0800 ;
        RECT 1.3800 1.8000 1.4700 2.0800 ;
        RECT 1.9000 1.8000 1.9900 2.0800 ;
        RECT 2.4200 1.8000 2.5100 2.0800 ;
        RECT 2.9400 1.8000 3.0300 2.0800 ;
        RECT 3.4600 1.8000 3.5500 2.0800 ;
        RECT 3.9800 1.8000 4.0700 2.0800 ;
        RECT 4.5700 1.8000 4.6600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 4.8900 1.8300 8.1000 1.9200 ;
      RECT 8.0100 1.4850 8.1000 1.8300 ;
      RECT 0.0800 1.6200 4.9800 1.7100 ;
      RECT 4.8900 1.7100 4.9800 1.8300 ;
      RECT 4.8900 1.5500 4.9800 1.6200 ;
      RECT 5.4100 1.4850 5.5000 1.8300 ;
      RECT 5.9300 1.4850 6.0200 1.8300 ;
      RECT 6.4500 1.4850 6.5400 1.8300 ;
      RECT 6.9700 1.4850 7.0600 1.8300 ;
      RECT 7.4900 1.4850 7.5800 1.8300 ;
      RECT 0.0800 1.7100 0.1700 1.9900 ;
      RECT 0.6000 1.7100 0.6900 1.9900 ;
      RECT 1.1200 1.7100 1.2100 1.9900 ;
      RECT 1.6400 1.7100 1.7300 1.9900 ;
      RECT 2.1600 1.7100 2.2500 1.9900 ;
      RECT 2.6800 1.7100 2.7700 1.9900 ;
      RECT 3.2000 1.7100 3.2900 1.9900 ;
      RECT 3.7200 1.7100 3.8100 1.9900 ;
      RECT 4.2400 1.7100 4.3300 1.9900 ;
  END
END AOI32_X6M_A12TH

MACRO BENC_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 15.2450 2.7200 ;
        RECT 0.2800 2.0450 0.5000 2.0800 ;
        RECT 1.6750 2.0400 1.8450 2.0800 ;
        RECT 11.6250 2.0050 11.7550 2.0800 ;
        RECT 12.1550 1.7750 12.2550 2.0800 ;
        RECT 12.6750 1.7600 12.7750 2.0800 ;
        RECT 13.1950 1.7600 13.2950 2.0800 ;
        RECT 13.7150 1.7600 13.8150 2.0800 ;
        RECT 14.2350 1.7600 14.3350 2.0800 ;
        RECT 14.7550 1.7600 14.8550 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 15.2450 0.3200 ;
        RECT 6.4250 0.3200 6.6350 0.3550 ;
        RECT 6.9450 0.3200 7.1550 0.3550 ;
        RECT 10.0150 0.3200 10.2250 0.3500 ;
        RECT 10.5200 0.3200 10.7300 0.3500 ;
        RECT 11.6150 0.3200 11.7550 0.5550 ;
        RECT 12.1550 0.3200 12.2550 0.6450 ;
        RECT 12.6400 0.3200 12.8100 0.5200 ;
        RECT 13.1600 0.3200 13.3300 0.5200 ;
        RECT 13.6800 0.3200 13.8500 0.5200 ;
        RECT 14.2000 0.3200 14.3700 0.5200 ;
        RECT 14.7200 0.3200 14.8900 0.5200 ;
    END
  END VSS

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.1450 0.3500 1.6500 ;
        RECT 0.2400 1.6500 5.7900 1.7400 ;
        RECT 5.6900 1.0500 5.7900 1.6500 ;
        RECT 5.6900 0.9500 6.0200 1.0500 ;
    END
    ANTENNAGATEAREA 0.1644 ;
  END M0

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.6200 0.8500 9.7800 1.2300 ;
        RECT 7.2100 1.2300 9.9100 1.3900 ;
        RECT 7.2100 0.6800 9.9100 0.8500 ;
        RECT 7.2100 1.3900 7.3300 1.5600 ;
        RECT 7.7300 1.3900 7.8300 1.5600 ;
        RECT 8.2500 1.3900 8.3500 1.5600 ;
        RECT 8.7700 1.3900 8.8700 1.5600 ;
        RECT 9.2900 1.3900 9.3900 1.5600 ;
        RECT 9.8000 1.3900 9.9100 1.5600 ;
    END
    ANTENNADIFFAREA 1.84135 ;
  END AN

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.4150 1.2250 15.1150 1.3850 ;
        RECT 12.4150 1.3850 12.5150 1.7200 ;
        RECT 12.9350 1.3850 13.0350 1.7200 ;
        RECT 13.4550 1.3850 13.5550 1.7200 ;
        RECT 13.9750 1.3850 14.0750 1.7200 ;
        RECT 14.4950 1.3850 14.5950 1.7200 ;
        RECT 15.0150 1.3850 15.1150 1.7200 ;
        RECT 14.9550 0.8700 15.1150 1.2250 ;
        RECT 12.4150 0.7100 15.1150 0.8700 ;
        RECT 12.9350 0.4550 13.0350 0.7100 ;
        RECT 13.4550 0.4550 13.5550 0.7100 ;
        RECT 12.4150 0.4500 12.5150 0.7100 ;
        RECT 13.9750 0.4500 14.0750 0.7100 ;
        RECT 14.4950 0.4500 14.5950 0.7100 ;
        RECT 15.0150 0.4500 15.1150 0.7100 ;
    END
    ANTENNADIFFAREA 1.885 ;
  END SN

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.5300 1.2500 11.1050 1.3500 ;
        RECT 10.5300 1.1000 10.6300 1.2500 ;
        RECT 11.0050 0.9100 11.1050 1.2500 ;
        RECT 10.2150 1.0000 10.6300 1.1000 ;
    END
    ANTENNAGATEAREA 0.0993 ;
  END M2

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7350 1.2100 1.9500 1.3100 ;
        RECT 1.8400 1.3100 1.9500 1.4700 ;
        RECT 1.7350 1.0350 1.8450 1.2100 ;
        RECT 1.8400 1.4700 5.5900 1.5600 ;
        RECT 5.4900 1.1500 5.5900 1.4700 ;
        RECT 5.4100 1.0500 5.5900 1.1500 ;
    END
    ANTENNAGATEAREA 0.2085 ;
  END M1

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8200 0.8300 4.9800 1.2200 ;
        RECT 2.6050 1.2200 4.9800 1.2400 ;
        RECT 2.6050 0.6700 5.3650 0.8300 ;
        RECT 2.6050 1.2400 5.3950 1.3800 ;
    END
    ANTENNADIFFAREA 1.878625 ;
  END X2
  OBS
    LAYER M1 ;
      RECT 0.5400 1.4400 0.7550 1.5550 ;
      RECT 0.6600 0.7900 0.7550 1.4400 ;
      RECT 0.5500 0.6700 0.7550 0.7900 ;
      RECT 1.5550 0.8400 2.0650 0.9300 ;
      RECT 1.9650 0.9300 2.0650 1.0050 ;
      RECT 1.9650 1.0050 2.3350 1.0950 ;
      RECT 0.8450 1.4650 1.6450 1.5550 ;
      RECT 1.5550 0.9300 1.6450 1.4650 ;
      RECT 0.8450 0.7900 0.9450 1.4650 ;
      RECT 0.8450 0.6700 1.0500 0.7900 ;
      RECT 2.4250 0.9900 4.4000 1.0800 ;
      RECT 2.0650 1.2550 2.5150 1.3450 ;
      RECT 2.4250 1.0800 2.5150 1.2550 ;
      RECT 2.4250 0.7500 2.5150 0.9900 ;
      RECT 2.0650 0.6600 2.5150 0.7500 ;
      RECT 5.4550 0.6600 6.1450 0.7700 ;
      RECT 6.0650 1.4550 6.1950 1.5550 ;
      RECT 6.0650 1.3550 6.4950 1.4550 ;
      RECT 6.4000 1.2100 6.4950 1.3550 ;
      RECT 6.4000 1.0400 6.9300 1.2100 ;
      RECT 6.4000 0.7700 6.4950 1.0400 ;
      RECT 6.2350 0.6600 6.4950 0.7700 ;
      RECT 7.0200 0.9950 9.2500 1.0850 ;
      RECT 6.6700 1.4450 7.1200 1.5450 ;
      RECT 7.0200 1.0850 7.1200 1.4450 ;
      RECT 7.0200 0.7950 7.1200 0.9950 ;
      RECT 6.6800 0.6950 7.1200 0.7950 ;
      RECT 10.0150 1.3400 10.4300 1.4400 ;
      RECT 10.3000 1.4400 10.4300 1.5350 ;
      RECT 10.0150 0.8100 10.4450 0.9100 ;
      RECT 10.3150 0.7050 10.4450 0.8100 ;
      RECT 5.8800 1.6500 10.1050 1.7400 ;
      RECT 10.0150 1.4400 10.1050 1.6500 ;
      RECT 10.0150 0.9100 10.1050 1.3400 ;
      RECT 5.8800 1.2550 5.9700 1.6500 ;
      RECT 5.8800 1.1550 6.2650 1.2550 ;
      RECT 6.1650 0.9100 6.2650 1.1550 ;
      RECT 1.3650 0.4800 10.6800 0.5700 ;
      RECT 10.5800 0.5700 10.6800 0.7550 ;
      RECT 10.5800 0.7550 10.8300 0.8550 ;
      RECT 10.7300 0.8550 10.8300 1.1200 ;
      RECT 1.2750 1.2650 1.4650 1.3750 ;
      RECT 1.3650 1.1500 1.4650 1.2650 ;
      RECT 1.0850 1.0500 1.4650 1.1500 ;
      RECT 1.3650 0.5700 1.4650 1.0500 ;
      RECT 10.7800 0.4800 11.5100 0.5800 ;
      RECT 11.3000 0.4700 11.5100 0.4800 ;
      RECT 11.3150 1.9200 11.5300 1.9300 ;
      RECT 10.5250 1.8200 11.5300 1.9200 ;
      RECT 10.8000 1.4600 11.3900 1.5500 ;
      RECT 11.2900 1.0500 11.3900 1.4600 ;
      RECT 11.2900 0.9500 11.5450 1.0500 ;
      RECT 0.0450 0.9900 0.1350 1.8300 ;
      RECT 0.0450 0.5800 0.1900 0.8900 ;
      RECT 0.0450 0.8900 0.5650 0.9900 ;
      RECT 0.4650 0.9900 0.5650 1.1000 ;
      RECT 0.0450 0.4800 1.2400 0.5800 ;
      RECT 1.1400 0.5800 1.2400 0.6700 ;
      RECT 0.0450 1.8300 10.4150 1.9200 ;
      RECT 10.3150 1.7300 10.4150 1.8300 ;
      RECT 10.3150 1.6400 10.9050 1.7300 ;
      RECT 10.8000 1.5500 10.9050 1.6400 ;
      RECT 11.0400 1.6400 11.7500 1.7300 ;
      RECT 11.6500 1.1850 11.7500 1.6400 ;
      RECT 11.6500 1.0850 12.0150 1.1850 ;
      RECT 11.6500 0.7850 11.7500 1.0850 ;
      RECT 11.0400 0.6850 11.7500 0.7850 ;
      RECT 12.1350 0.9850 14.4500 1.0850 ;
      RECT 11.8950 1.4800 11.9950 1.8250 ;
      RECT 11.8750 0.4650 12.0150 0.7600 ;
      RECT 11.8950 1.3800 12.2350 1.4800 ;
      RECT 12.1350 1.0850 12.2350 1.3800 ;
      RECT 12.1350 0.8600 12.2350 0.9850 ;
      RECT 11.8750 0.7600 12.2350 0.8600 ;
  END
END BENC_X11M_A12TH

MACRO BENC_X16M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 21.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 21.6450 2.7200 ;
        RECT 7.2700 2.0600 7.4800 2.0800 ;
        RECT 13.9250 2.0450 14.1450 2.0800 ;
        RECT 2.3400 2.0400 2.5600 2.0800 ;
        RECT 2.8700 2.0400 3.0800 2.0800 ;
        RECT 3.3900 2.0400 3.6000 2.0800 ;
        RECT 3.9100 2.0400 4.1200 2.0800 ;
        RECT 4.4300 2.0400 4.6400 2.0800 ;
        RECT 4.9500 2.0400 5.1600 2.0800 ;
        RECT 5.4700 2.0400 5.6800 2.0800 ;
        RECT 5.9900 2.0400 6.2000 2.0800 ;
        RECT 6.5100 2.0400 6.7200 2.0800 ;
        RECT 9.7700 2.0100 9.9800 2.0800 ;
        RECT 9.2700 1.9150 9.4400 2.0800 ;
        RECT 15.7100 1.8200 15.8000 2.0800 ;
        RECT 17.7800 1.7600 17.8800 2.0800 ;
        RECT 18.3000 1.7600 18.4000 2.0800 ;
        RECT 18.8200 1.7600 18.9200 2.0800 ;
        RECT 19.3400 1.7600 19.4400 2.0800 ;
        RECT 19.8600 1.7600 19.9600 2.0800 ;
        RECT 20.3800 1.7600 20.4800 2.0800 ;
        RECT 20.9000 1.7600 21.0000 2.0800 ;
        RECT 21.4200 1.7600 21.5200 2.0800 ;
        RECT 14.6450 1.7550 14.7350 2.0800 ;
        RECT 16.7400 1.6700 16.8600 2.0800 ;
        RECT 17.2600 1.6100 17.3600 2.0800 ;
        RECT 16.2700 1.6050 16.3700 2.0800 ;
    END
  END VDD

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.3750 0.9100 13.6250 1.2300 ;
        RECT 10.0850 1.2300 13.6250 1.2850 ;
        RECT 10.0850 0.6800 13.8250 0.9100 ;
        RECT 10.0850 1.2850 13.8250 1.4800 ;
    END
    ANTENNADIFFAREA 2.6 ;
  END AN

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 15.3650 1.2500 15.9150 1.3500 ;
        RECT 15.8150 1.0750 15.9150 1.2500 ;
        RECT 15.3650 0.9400 15.4650 1.2500 ;
        RECT 15.8150 0.9750 16.1750 1.0750 ;
        RECT 14.9650 0.8400 15.4650 0.9400 ;
        RECT 14.9650 0.9400 15.0650 1.2350 ;
        RECT 14.4650 1.2350 15.0650 1.3350 ;
        RECT 14.4650 1.0800 14.5650 1.2350 ;
        RECT 14.1250 0.9800 14.5650 1.0800 ;
    END
    ANTENNAGATEAREA 0.177 ;
  END M2

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5850 0.9300 6.7900 1.1900 ;
        RECT 6.5850 1.1900 6.6850 1.4700 ;
        RECT 0.8300 1.4700 6.6850 1.5600 ;
        RECT 1.2500 1.4050 1.4200 1.4700 ;
        RECT 0.8300 0.8450 0.9400 1.4700 ;
    END
    ANTENNAGATEAREA 0.3369 ;
  END M1

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 21.0050 0.8200 21.2550 1.2950 ;
        RECT 17.4850 1.2950 21.2550 1.6050 ;
        RECT 17.4650 0.5100 21.2550 0.8200 ;
        RECT 21.1000 1.6050 21.2550 1.6850 ;
    END
    ANTENNADIFFAREA 2.6 ;
  END SN

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5750 0.9750 6.4400 1.1800 ;
        RECT 2.6300 1.1800 6.4400 1.2250 ;
        RECT 4.5750 0.8400 4.8550 0.9750 ;
        RECT 5.2300 0.6600 5.3850 0.9750 ;
        RECT 5.7450 0.6600 5.9100 0.9750 ;
        RECT 6.2750 0.6600 6.4400 0.9750 ;
        RECT 2.6300 1.2250 4.8900 1.3800 ;
        RECT 5.2300 1.2250 5.4000 1.3800 ;
        RECT 5.7500 1.2250 5.9200 1.3800 ;
        RECT 6.2700 1.2250 6.4400 1.3800 ;
        RECT 2.6100 0.6800 4.8550 0.8400 ;
    END
    ANTENNADIFFAREA 2.6 ;
  END X2

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 1.2900 0.4250 1.3900 ;
        RECT 0.3350 1.3900 0.4250 1.6500 ;
        RECT 0.2350 1.0350 0.3500 1.2900 ;
        RECT 0.3350 1.6500 7.4150 1.7400 ;
        RECT 7.2750 1.5600 7.4150 1.6500 ;
        RECT 7.2750 1.4700 8.4250 1.5600 ;
        RECT 8.3350 1.1500 8.4250 1.4700 ;
        RECT 7.6850 1.0500 8.4250 1.1500 ;
    END
    ANTENNAGATEAREA 0.267 ;
  END M0

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 21.6450 0.3200 ;
        RECT 0.2900 0.3200 0.5000 0.3800 ;
        RECT 1.7950 0.3200 2.0400 0.3800 ;
        RECT 2.3300 0.3200 2.5750 0.3800 ;
        RECT 7.2700 0.3200 7.4800 0.3550 ;
        RECT 7.7900 0.3200 8.0000 0.3550 ;
        RECT 16.7400 0.3200 16.8400 0.6400 ;
        RECT 17.2550 0.3200 17.3550 0.6400 ;
        RECT 21.4150 0.3200 21.5150 0.6400 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.5800 1.3300 0.7350 1.5550 ;
      RECT 0.6450 0.7500 0.7350 1.3300 ;
      RECT 0.5300 0.6600 0.7350 0.7500 ;
      RECT 1.0400 1.2050 1.1500 1.3800 ;
      RECT 1.0400 1.1300 1.4800 1.2050 ;
      RECT 1.0400 1.1150 2.2850 1.1300 ;
      RECT 1.3850 1.0300 2.2850 1.1150 ;
      RECT 1.0400 0.7550 1.1300 1.1150 ;
      RECT 0.8750 0.6600 1.1300 0.7550 ;
      RECT 2.3950 0.9900 4.1600 1.0800 ;
      RECT 1.5300 1.2800 2.4850 1.3700 ;
      RECT 2.3950 1.0800 2.4850 1.2800 ;
      RECT 2.3950 0.8800 2.4850 0.9900 ;
      RECT 1.5250 0.7900 2.4850 0.8800 ;
      RECT 7.0650 1.2700 8.2400 1.3800 ;
      RECT 7.0650 1.3800 7.1650 1.4850 ;
      RECT 7.0700 0.7500 7.1900 0.8350 ;
      RECT 7.0700 0.6800 8.9100 0.7500 ;
      RECT 8.6700 0.7500 8.9100 0.7700 ;
      RECT 7.0700 0.6600 8.7600 0.6800 ;
      RECT 7.7300 1.6500 8.6850 1.7400 ;
      RECT 8.5800 1.4850 8.6850 1.6500 ;
      RECT 8.5150 1.3850 8.6850 1.4850 ;
      RECT 8.5150 0.9900 8.6100 1.3850 ;
      RECT 8.5150 0.9650 9.7100 0.9900 ;
      RECT 9.0450 0.9900 9.7100 1.0650 ;
      RECT 8.5150 0.9500 9.1450 0.9650 ;
      RECT 8.4000 0.8800 9.1450 0.9500 ;
      RECT 8.4000 0.8400 8.6100 0.8800 ;
      RECT 9.8750 1.0200 12.9250 1.1200 ;
      RECT 9.0050 1.3350 9.9750 1.4350 ;
      RECT 9.8750 1.1200 9.9750 1.3350 ;
      RECT 9.8750 0.7700 9.9750 1.0200 ;
      RECT 9.0100 0.6800 9.9750 0.7700 ;
      RECT 13.9250 1.2150 14.3400 1.3150 ;
      RECT 14.2500 1.3150 14.3400 1.6900 ;
      RECT 13.9250 0.6900 14.3400 0.8750 ;
      RECT 9.7900 1.6400 14.0150 1.7300 ;
      RECT 13.9250 1.3150 14.0150 1.6400 ;
      RECT 13.9250 0.8750 14.0150 1.2150 ;
      RECT 9.7900 1.6350 9.8800 1.6400 ;
      RECT 8.8150 1.5450 9.8800 1.6350 ;
      RECT 8.8150 1.1900 8.9150 1.5450 ;
      RECT 8.7100 1.0800 8.9150 1.1900 ;
      RECT 14.4400 1.4400 15.2750 1.5300 ;
      RECT 15.1850 1.0500 15.2750 1.4400 ;
      RECT 0.0550 1.8300 9.0800 1.9200 ;
      RECT 8.9800 1.8150 9.0800 1.8300 ;
      RECT 8.9800 1.7250 9.6800 1.8150 ;
      RECT 9.5900 1.8150 9.6800 1.8300 ;
      RECT 0.0550 0.9350 0.1450 1.5450 ;
      RECT 0.0550 0.5700 0.1900 0.8400 ;
      RECT 0.0550 1.5450 0.2350 1.8300 ;
      RECT 0.0550 0.8400 0.5400 0.9350 ;
      RECT 0.4500 0.9350 0.5400 1.0500 ;
      RECT 0.0550 0.5200 1.0700 0.5700 ;
      RECT 0.0550 0.4800 1.3850 0.5200 ;
      RECT 0.9800 0.4300 1.3850 0.4800 ;
      RECT 9.5900 1.8300 14.5300 1.9200 ;
      RECT 14.4400 1.5300 14.5300 1.8300 ;
      RECT 14.4300 0.6600 15.6450 0.7500 ;
      RECT 15.5550 0.7500 15.6450 1.1200 ;
      RECT 6.8000 1.3200 6.9700 1.5200 ;
      RECT 6.8800 0.8200 6.9700 1.3200 ;
      RECT 6.7900 0.5700 6.9700 0.8200 ;
      RECT 2.3800 0.5700 2.4750 0.6100 ;
      RECT 1.2200 0.6100 2.4750 0.7000 ;
      RECT 1.2200 0.7000 1.3100 0.9800 ;
      RECT 2.3800 0.4800 14.5200 0.5700 ;
      RECT 14.4300 0.5700 14.5200 0.6600 ;
      RECT 14.7500 0.7500 14.8400 1.1400 ;
      RECT 15.7550 0.5700 15.8450 0.8300 ;
      RECT 14.6100 0.4800 16.4250 0.5700 ;
      RECT 14.6100 0.4100 14.7950 0.4800 ;
      RECT 16.2650 0.9600 17.1500 1.0600 ;
      RECT 15.1500 1.6400 16.1100 1.7300 ;
      RECT 16.0100 1.3150 16.1100 1.6400 ;
      RECT 16.0100 1.2250 16.3650 1.3150 ;
      RECT 16.2650 1.0600 16.3650 1.2250 ;
      RECT 16.2650 0.7900 16.3650 0.9600 ;
      RECT 15.9400 0.6900 16.3650 0.7900 ;
      RECT 15.1500 1.7300 15.3200 1.9300 ;
      RECT 17.2550 1.0300 20.3850 1.1200 ;
      RECT 16.4800 1.2800 17.3550 1.3800 ;
      RECT 17.2550 1.1200 17.3550 1.2800 ;
      RECT 17.2550 0.8500 17.3550 1.0300 ;
      RECT 16.4800 0.7500 17.3550 0.8500 ;
      RECT 16.4800 1.3800 16.5800 1.5450 ;
      RECT 16.4800 0.6600 16.5800 0.7500 ;
      RECT 17.0000 1.3800 17.1000 1.7550 ;
      RECT 17.0000 0.4500 17.1000 0.7500 ;
  END
END BENC_X16M_A12TH

MACRO BENC_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 5.5050 1.8300 5.6050 2.0800 ;
        RECT 6.0250 1.7500 6.1250 2.0800 ;
    END
  END VDD

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 1.0100 4.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.105 ;
  END M2

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.6500 1.1900 ;
        RECT 1.4500 0.8500 1.7900 0.9500 ;
        RECT 1.6900 0.7500 1.7900 0.8500 ;
        RECT 1.6900 0.6600 2.7050 0.7500 ;
        RECT 2.5900 0.7500 2.7050 1.1650 ;
    END
    ANTENNAGATEAREA 0.2187 ;
  END M1

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0500 0.9500 6.1500 1.2500 ;
        RECT 5.7650 1.2500 6.1500 1.3500 ;
        RECT 5.7600 0.8500 6.1500 0.9500 ;
        RECT 5.7650 1.3500 5.8650 1.7400 ;
        RECT 5.7600 0.4400 5.8600 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END AN

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.2500 ;
        RECT 2.0150 1.2500 2.3500 1.3500 ;
        RECT 1.9500 0.8400 2.3500 0.9500 ;
        RECT 2.0150 1.3500 2.1150 1.5500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END X2

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6500 0.8100 4.1500 0.9500 ;
        RECT 4.0500 0.9500 4.1500 1.2500 ;
        RECT 3.7150 1.2500 4.1500 1.3500 ;
        RECT 3.7150 1.3500 3.8150 1.5600 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END SN

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 1.4500 2.9450 1.5500 ;
        RECT 2.2250 1.5500 2.3350 1.6400 ;
        RECT 2.8050 0.9250 2.9450 1.4500 ;
        RECT 0.3700 1.6400 2.3350 1.7400 ;
        RECT 0.3700 1.3600 0.4700 1.6400 ;
        RECT 0.2350 1.2600 0.4700 1.3600 ;
        RECT 0.2350 1.0400 0.3350 1.2600 ;
    END
    ANTENNAGATEAREA 0.1776 ;
  END M0

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.2850 0.3200 0.4950 0.3900 ;
        RECT 1.6450 0.3200 1.8550 0.3500 ;
        RECT 2.2450 0.3200 2.6150 0.3650 ;
        RECT 6.0250 0.3200 6.1250 0.6400 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.5900 1.3500 0.7000 1.5500 ;
      RECT 0.5900 1.2600 0.9000 1.3500 ;
      RECT 0.8100 0.9750 0.9000 1.2600 ;
      RECT 0.6450 0.8850 0.9000 0.9750 ;
      RECT 0.6450 0.7500 0.7350 0.8850 ;
      RECT 0.5350 0.6600 0.7350 0.7500 ;
      RECT 1.7650 1.0650 2.0350 1.1550 ;
      RECT 0.8050 1.4600 1.8650 1.5500 ;
      RECT 1.7650 1.1550 1.8650 1.4600 ;
      RECT 0.8050 1.4400 1.1250 1.4600 ;
      RECT 1.0350 0.7700 1.1250 1.4400 ;
      RECT 0.8250 0.6600 1.1250 0.7700 ;
      RECT 2.4450 1.6400 3.1700 1.7400 ;
      RECT 3.4000 1.0450 3.8500 1.1450 ;
      RECT 3.2350 1.2600 3.5000 1.3700 ;
      RECT 3.4000 1.1450 3.5000 1.2600 ;
      RECT 3.4000 0.7600 3.5000 1.0450 ;
      RECT 2.9300 0.6600 3.5000 0.7600 ;
      RECT 3.3550 1.6500 4.1100 1.7400 ;
      RECT 4.0200 1.5600 4.1100 1.6500 ;
      RECT 4.0200 1.4700 4.3300 1.5600 ;
      RECT 4.2400 0.7200 4.3300 1.4700 ;
      RECT 3.3550 1.5500 3.4450 1.6500 ;
      RECT 3.0400 1.4600 3.4450 1.5500 ;
      RECT 3.0400 1.0850 3.1300 1.4600 ;
      RECT 3.0400 0.9850 3.2700 1.0850 ;
      RECT 4.2100 1.6500 4.5550 1.7400 ;
      RECT 4.4550 1.3700 4.5550 1.6500 ;
      RECT 4.4550 1.2800 5.0350 1.3700 ;
      RECT 4.9350 0.9150 5.0350 1.2800 ;
      RECT 0.0550 1.8300 4.3100 1.9200 ;
      RECT 4.2100 1.7400 4.3100 1.8300 ;
      RECT 0.0550 1.4700 0.1950 1.8300 ;
      RECT 0.0550 0.9300 0.1450 1.4700 ;
      RECT 0.0550 0.5700 0.1950 0.8400 ;
      RECT 0.0550 0.8400 0.5350 0.9300 ;
      RECT 0.4350 0.9300 0.5350 1.0700 ;
      RECT 0.4350 1.0700 0.6600 1.1700 ;
      RECT 0.0550 0.4800 1.2550 0.5700 ;
      RECT 1.3900 0.4800 4.5750 0.5700 ;
      RECT 4.4750 0.5700 4.5750 0.6600 ;
      RECT 4.4750 0.6600 5.2600 0.7600 ;
      RECT 5.1600 0.7600 5.2600 1.1150 ;
      RECT 1.2250 0.7500 1.3150 1.2800 ;
      RECT 1.2250 1.2800 1.5600 1.3700 ;
      RECT 1.2250 0.6600 1.4900 0.7500 ;
      RECT 1.3900 0.5700 1.4900 0.6600 ;
      RECT 4.6900 1.4600 5.3650 1.5600 ;
      RECT 5.2650 1.3100 5.3650 1.4600 ;
      RECT 5.5000 1.0500 5.9250 1.1500 ;
      RECT 4.9300 1.6500 5.5900 1.7400 ;
      RECT 5.5000 1.1500 5.5900 1.6500 ;
      RECT 5.5000 0.5700 5.5900 1.0500 ;
      RECT 4.6750 0.4800 5.5900 0.5700 ;
      RECT 4.4300 1.8300 5.0200 1.9200 ;
      RECT 4.9300 1.7400 5.0200 1.8300 ;
      RECT 4.6750 0.4600 4.9100 0.4800 ;
  END
END BENC_X2M_A12TH

MACRO BENC_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.2450 2.7200 ;
        RECT 2.4050 2.0200 2.6150 2.0800 ;
        RECT 2.9450 2.0200 3.3150 2.0800 ;
        RECT 7.2350 1.9900 7.3350 2.0800 ;
        RECT 7.7550 1.7600 7.8550 2.0800 ;
        RECT 6.2050 1.7550 6.3050 2.0800 ;
        RECT 6.7350 1.7150 6.8350 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.2450 0.3200 ;
        RECT 1.6400 0.3200 1.8100 0.3900 ;
        RECT 4.4550 0.3200 4.6800 0.3900 ;
        RECT 5.9000 0.3200 6.0900 0.3900 ;
        RECT 7.2350 0.3200 7.3350 0.4100 ;
        RECT 7.7550 0.3200 7.8550 0.6400 ;
    END
  END VSS

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.2500 3.6650 1.3500 ;
        RECT 3.2500 1.3500 3.3500 1.6500 ;
        RECT 3.5650 0.9100 3.6650 1.2500 ;
        RECT 0.3350 1.6500 3.3500 1.7400 ;
        RECT 0.3350 1.3900 0.4250 1.6500 ;
        RECT 0.2300 1.3000 0.4250 1.3900 ;
        RECT 0.2300 1.1300 0.3500 1.3000 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END M0

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2000 0.8500 2.8600 0.9500 ;
        RECT 2.7600 0.9500 2.8600 1.2500 ;
        RECT 2.2000 0.7000 2.3000 0.8500 ;
        RECT 2.7200 0.7000 2.8600 0.8500 ;
        RECT 2.1650 1.2500 2.8600 1.3800 ;
    END
    ANTENNADIFFAREA 0.59865 ;
  END X2

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4950 1.2500 8.1150 1.3500 ;
        RECT 7.4950 1.3500 7.5950 1.7450 ;
        RECT 8.0150 1.3500 8.1150 1.7450 ;
        RECT 8.0150 0.9500 8.1150 1.2500 ;
        RECT 7.4900 0.8500 8.1150 0.9500 ;
        RECT 7.4900 0.4500 7.5900 0.8500 ;
        RECT 8.0150 0.4500 8.1150 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END SN

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 1.0500 3.4250 1.1500 ;
        RECT 3.0500 1.1500 3.1500 1.4700 ;
        RECT 3.3250 0.9050 3.4250 1.0500 ;
        RECT 1.6500 1.4700 3.1500 1.5600 ;
        RECT 1.6500 1.3200 1.7500 1.4700 ;
        RECT 1.5600 1.2100 1.7500 1.3200 ;
        RECT 1.5600 1.0300 1.6750 1.2100 ;
    END
    ANTENNAGATEAREA 0.1089 ;
  END M1

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0100 1.0500 6.5450 1.1500 ;
    END
    ANTENNAGATEAREA 0.06 ;
  END M2

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7750 1.2500 5.4000 1.3500 ;
        RECT 4.7750 1.3500 4.8750 1.4900 ;
        RECT 5.2900 1.3500 5.4000 1.4900 ;
        RECT 5.3000 0.9500 5.4000 1.2500 ;
        RECT 4.7800 0.8500 5.4000 0.9500 ;
        RECT 4.7800 0.7050 4.8800 0.8500 ;
        RECT 5.3000 0.7050 5.4000 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END AN
  OBS
    LAYER M1 ;
      RECT 0.5450 1.4200 0.7850 1.5350 ;
      RECT 0.6950 0.7900 0.7850 1.4200 ;
      RECT 0.5650 0.6800 0.7850 0.7900 ;
      RECT 1.3800 0.8500 1.8850 0.9400 ;
      RECT 1.7750 0.9400 1.8850 1.1000 ;
      RECT 0.8750 1.4700 1.4700 1.5600 ;
      RECT 1.3800 0.9400 1.4700 1.4700 ;
      RECT 0.8750 0.6600 0.9950 1.4700 ;
      RECT 1.9750 1.0500 2.6500 1.1500 ;
      RECT 1.8850 1.2800 2.0750 1.3800 ;
      RECT 1.9750 1.1500 2.0750 1.2800 ;
      RECT 1.9750 0.7500 2.0750 1.0500 ;
      RECT 1.8700 0.6600 2.0750 0.7500 ;
      RECT 3.1550 0.6600 3.9050 0.7500 ;
      RECT 3.7550 0.9700 3.8550 1.4450 ;
      RECT 3.7550 0.8800 4.4500 0.9700 ;
      RECT 4.3600 0.9700 4.4500 1.1850 ;
      RECT 4.0200 0.6800 4.1200 0.8800 ;
      RECT 4.5750 1.0450 5.1100 1.1450 ;
      RECT 4.2150 1.3800 4.6650 1.4900 ;
      RECT 4.5750 1.1450 4.6650 1.3800 ;
      RECT 4.5750 0.7500 4.6650 1.0450 ;
      RECT 4.2150 0.6600 4.6650 0.7500 ;
      RECT 4.2150 0.7500 4.4050 0.7700 ;
      RECT 0.0500 1.8900 5.9450 1.9200 ;
      RECT 5.6600 1.9200 5.9450 1.9900 ;
      RECT 0.0500 1.8300 5.7600 1.8900 ;
      RECT 0.0500 1.5450 0.1700 1.8300 ;
      RECT 0.0500 1.0050 0.1400 1.5450 ;
      RECT 0.0500 0.5700 0.1750 0.9050 ;
      RECT 1.0900 1.9200 1.2900 1.9800 ;
      RECT 0.0500 0.9050 0.5950 1.0050 ;
      RECT 0.0500 0.4800 1.2950 0.5700 ;
      RECT 0.8750 0.4600 1.2950 0.4800 ;
      RECT 5.4900 0.8600 6.2150 0.9500 ;
      RECT 1.4050 0.4800 5.5900 0.5700 ;
      RECT 5.4900 0.5700 5.5900 0.8600 ;
      RECT 1.0850 1.2700 1.2900 1.3800 ;
      RECT 1.0850 0.7600 1.1750 1.2700 ;
      RECT 1.0850 0.6600 1.5050 0.7600 ;
      RECT 1.4050 0.5700 1.5050 0.6600 ;
      RECT 5.6800 0.4800 6.3400 0.5800 ;
      RECT 5.6800 0.4100 5.7900 0.4800 ;
      RECT 5.4900 1.3100 6.7550 1.4100 ;
      RECT 6.6650 0.9200 6.7550 1.3100 ;
      RECT 6.4700 0.8300 6.7550 0.9200 ;
      RECT 6.4700 0.7050 6.5800 0.8300 ;
      RECT 3.9850 1.5800 5.5900 1.6700 ;
      RECT 5.4900 1.4100 5.5900 1.5800 ;
      RECT 3.9850 1.1700 4.0850 1.5800 ;
      RECT 3.9850 1.0600 4.1850 1.1700 ;
      RECT 5.6800 1.5150 6.9350 1.6050 ;
      RECT 6.8450 0.7200 6.9350 1.5150 ;
      RECT 6.7300 0.6300 6.9350 0.7200 ;
      RECT 6.7300 0.5500 6.8300 0.6300 ;
      RECT 6.4300 0.4600 6.8300 0.5500 ;
      RECT 5.6800 1.6050 5.7700 1.7200 ;
      RECT 6.4650 1.6050 6.5650 1.9150 ;
      RECT 7.0500 1.0500 7.9050 1.1500 ;
      RECT 6.9550 1.7050 7.1400 1.8050 ;
      RECT 7.0500 1.1500 7.1400 1.7050 ;
      RECT 7.0500 0.5300 7.1400 1.0500 ;
      RECT 6.9600 0.4400 7.1400 0.5300 ;
  END
END BENC_X3M_A12TH

MACRO BENC_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.8450 2.7200 ;
        RECT 2.1200 2.0200 2.3300 2.0800 ;
        RECT 2.6400 2.0200 2.8500 2.0800 ;
        RECT 3.1800 2.0200 3.5500 2.0800 ;
        RECT 7.5850 1.9900 7.6850 2.0800 ;
        RECT 7.0850 1.8950 7.1850 2.0800 ;
        RECT 8.1050 1.7600 8.2050 2.0800 ;
        RECT 8.6250 1.7600 8.7250 2.0800 ;
        RECT 6.5550 1.7500 6.6550 2.0800 ;
    END
  END VDD

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0100 1.2500 5.6350 1.3500 ;
        RECT 5.0100 1.3500 5.1100 1.4900 ;
        RECT 5.5300 1.3500 5.6350 1.4900 ;
        RECT 5.5350 0.9500 5.6350 1.2500 ;
        RECT 5.0150 0.8500 5.6350 0.9500 ;
        RECT 5.0150 0.6950 5.1150 0.8500 ;
        RECT 5.5350 0.6950 5.6350 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END AN

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.3650 1.0500 6.8950 1.1500 ;
    END
    ANTENNAGATEAREA 0.0684 ;
  END M2

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.0500 3.6600 1.1500 ;
        RECT 3.2500 1.1500 3.3500 1.4700 ;
        RECT 3.5600 0.9050 3.6600 1.0500 ;
        RECT 1.5900 1.4700 3.3500 1.5600 ;
        RECT 1.5900 1.0300 1.6900 1.4700 ;
    END
    ANTENNAGATEAREA 0.1275 ;
  END M1

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8450 1.2500 8.4650 1.3500 ;
        RECT 7.8450 1.3500 7.9450 1.7350 ;
        RECT 8.3650 1.3500 8.4650 1.7350 ;
        RECT 8.3650 0.9500 8.4650 1.2500 ;
        RECT 7.8400 0.8500 8.4650 0.9500 ;
        RECT 7.8400 0.4500 7.9400 0.8500 ;
        RECT 8.3650 0.4500 8.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END SN

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4350 0.8500 3.0950 0.9500 ;
        RECT 2.9950 0.9500 3.0950 1.2500 ;
        RECT 2.9550 0.6900 3.0950 0.8500 ;
        RECT 2.4350 0.6850 2.5350 0.8500 ;
        RECT 2.3700 1.2500 3.0950 1.3800 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END X2

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.2500 3.9500 1.3500 ;
        RECT 3.4500 1.3500 3.5500 1.6500 ;
        RECT 3.8400 0.9100 3.9500 1.2500 ;
        RECT 0.3350 1.6500 3.5500 1.7400 ;
        RECT 0.3350 1.3900 0.4250 1.6500 ;
        RECT 0.2300 1.3000 0.4250 1.3900 ;
        RECT 0.2300 1.1300 0.3500 1.3000 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END M0

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.8450 0.3200 ;
        RECT 1.6200 0.3200 1.8300 0.3750 ;
        RECT 6.2300 0.3200 6.4400 0.3550 ;
        RECT 7.0300 0.3200 7.2400 0.3300 ;
        RECT 7.5850 0.3200 7.6850 0.4100 ;
        RECT 8.1050 0.3200 8.2050 0.6400 ;
        RECT 8.6250 0.3200 8.7250 0.6400 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.5450 1.4200 0.7850 1.5350 ;
      RECT 0.6950 0.7900 0.7850 1.4200 ;
      RECT 0.5650 0.6800 0.7850 0.7900 ;
      RECT 1.3900 0.8500 1.9300 0.9400 ;
      RECT 1.8300 0.9400 1.9300 1.1750 ;
      RECT 0.8750 1.4700 1.4800 1.5600 ;
      RECT 1.3900 0.9400 1.4800 1.4700 ;
      RECT 0.8750 0.6600 0.9950 1.4700 ;
      RECT 2.1550 1.0500 2.8300 1.1500 ;
      RECT 1.8850 1.2800 2.2550 1.3800 ;
      RECT 2.1550 1.1500 2.2550 1.2800 ;
      RECT 2.1550 0.7500 2.2550 1.0500 ;
      RECT 1.8700 0.6600 2.2550 0.7500 ;
      RECT 3.3900 0.6600 4.1500 0.7500 ;
      RECT 3.9250 1.4500 4.1600 1.5500 ;
      RECT 4.0600 0.9300 4.1600 1.4500 ;
      RECT 4.0600 0.8400 4.6950 0.9300 ;
      RECT 4.6050 0.9300 4.6950 1.1850 ;
      RECT 4.2600 0.6600 4.3500 0.8400 ;
      RECT 4.8100 1.0450 5.3450 1.1450 ;
      RECT 4.4600 1.3800 4.9000 1.4900 ;
      RECT 4.8100 1.1450 4.9000 1.3800 ;
      RECT 4.8100 0.7500 4.9000 1.0450 ;
      RECT 4.4600 0.6600 4.9000 0.7500 ;
      RECT 0.0500 1.8900 6.2950 1.9200 ;
      RECT 6.0100 1.9200 6.2950 1.9900 ;
      RECT 0.0500 1.8300 6.1100 1.8900 ;
      RECT 0.0500 1.4800 0.2100 1.8300 ;
      RECT 0.0500 1.0050 0.1400 1.4800 ;
      RECT 0.0500 0.5700 0.1750 0.9050 ;
      RECT 1.0900 1.9200 1.2900 1.9800 ;
      RECT 0.0500 0.9050 0.5950 1.0050 ;
      RECT 0.0500 0.4800 1.2950 0.5700 ;
      RECT 0.8750 0.4600 1.2950 0.4800 ;
      RECT 5.7750 0.8600 6.5650 0.9500 ;
      RECT 1.4050 0.4800 5.8750 0.5700 ;
      RECT 5.7750 0.5700 5.8750 0.8600 ;
      RECT 1.0850 1.2700 1.3000 1.3800 ;
      RECT 1.0850 0.7600 1.1750 1.2700 ;
      RECT 1.0850 0.6600 1.5050 0.7600 ;
      RECT 1.4050 0.5700 1.5050 0.6600 ;
      RECT 5.9650 0.4800 6.6900 0.5800 ;
      RECT 5.7500 1.3100 7.1050 1.4100 ;
      RECT 7.0150 0.9200 7.1050 1.3100 ;
      RECT 6.8200 0.8300 7.1050 0.9200 ;
      RECT 6.8200 0.7050 6.9300 0.8300 ;
      RECT 4.2650 1.5800 5.8500 1.6700 ;
      RECT 5.7500 1.4100 5.8500 1.5800 ;
      RECT 4.2650 1.2150 4.3650 1.5800 ;
      RECT 4.2650 1.0200 4.3750 1.2150 ;
      RECT 5.9700 1.5150 7.2850 1.6050 ;
      RECT 7.1950 0.7200 7.2850 1.5150 ;
      RECT 7.0800 0.6300 7.2850 0.7200 ;
      RECT 7.0800 0.5700 7.1800 0.6300 ;
      RECT 6.7800 0.4800 7.1800 0.5700 ;
      RECT 6.8150 1.6050 6.9150 1.9150 ;
      RECT 7.4000 1.0500 8.2550 1.1500 ;
      RECT 7.3050 1.8200 7.4900 1.9200 ;
      RECT 7.4000 1.1500 7.4900 1.8200 ;
      RECT 7.4000 0.5300 7.4900 1.0500 ;
      RECT 7.3100 0.4400 7.4900 0.5300 ;
  END
END BENC_X4M_A12TH

MACRO BENC_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 11.0450 2.7200 ;
        RECT 0.2900 2.0450 0.5000 2.0800 ;
        RECT 2.3350 2.0400 2.5550 2.0800 ;
        RECT 8.7350 1.8400 8.8350 2.0800 ;
        RECT 8.2200 1.8300 8.3300 2.0800 ;
        RECT 9.2550 1.7600 9.3550 2.0800 ;
        RECT 9.7750 1.7600 9.8750 2.0800 ;
        RECT 10.2950 1.7600 10.3950 2.0800 ;
        RECT 10.8150 1.7600 10.9150 2.0800 ;
    END
  END VDD

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9850 1.5650 1.1900 ;
        RECT 1.4500 0.8950 2.0000 0.9850 ;
        RECT 1.9100 0.9850 2.0000 1.4700 ;
        RECT 1.9100 1.4700 4.3600 1.5600 ;
        RECT 4.2500 0.9550 4.3600 1.4700 ;
    END
    ANTENNAGATEAREA 0.1752 ;
  END M1

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.1550 0.4300 1.3900 ;
        RECT 0.3300 1.3900 0.4300 1.6500 ;
        RECT 0.3300 1.6500 4.5500 1.7400 ;
        RECT 4.4500 1.1700 4.5500 1.6500 ;
        RECT 4.4500 0.9450 4.6200 1.1700 ;
    END
    ANTENNAGATEAREA 0.1359 ;
  END M0

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8300 0.8000 3.9700 1.2400 ;
        RECT 2.6200 1.2400 3.9700 1.3800 ;
        RECT 2.6200 0.6600 3.9700 0.8000 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END X2

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9000 1.2500 7.1150 1.4050 ;
        RECT 6.9750 0.8200 7.1150 1.2500 ;
        RECT 5.9050 0.6800 7.1150 0.8200 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END AN

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5150 1.2400 10.7700 1.3800 ;
        RECT 9.5150 1.3800 9.6150 1.7350 ;
        RECT 10.0350 1.3800 10.1350 1.7350 ;
        RECT 10.5550 1.3800 10.6550 1.7350 ;
        RECT 10.6300 0.9600 10.7700 1.2400 ;
        RECT 9.5150 0.8200 10.7700 0.9600 ;
        RECT 10.0350 0.4400 10.1350 0.8200 ;
        RECT 10.5550 0.4400 10.6550 0.8200 ;
        RECT 9.5150 0.4300 9.6150 0.8200 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END SN

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.1950 1.0100 8.6950 1.1900 ;
    END
    ANTENNAGATEAREA 0.0852 ;
  END M2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 11.0450 0.3200 ;
        RECT 4.3650 0.3200 4.5750 0.3900 ;
        RECT 7.6800 0.3200 7.8300 0.4550 ;
        RECT 9.2550 0.3200 9.3550 0.7300 ;
        RECT 9.7750 0.3200 9.8750 0.6050 ;
        RECT 10.2950 0.3200 10.3950 0.6050 ;
        RECT 10.8150 0.3200 10.9150 0.6200 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.5550 1.4400 0.7650 1.5600 ;
      RECT 0.6650 0.7750 0.7650 1.4400 ;
      RECT 0.5600 0.6600 0.7650 0.7750 ;
      RECT 0.8800 1.4700 1.8200 1.5600 ;
      RECT 1.7100 1.0750 1.8200 1.4700 ;
      RECT 0.8800 0.6800 0.9750 1.4700 ;
      RECT 2.3500 0.9800 3.6950 1.0800 ;
      RECT 2.0900 1.2700 2.4500 1.3800 ;
      RECT 2.3500 1.0800 2.4500 1.2700 ;
      RECT 2.3500 0.7500 2.4500 0.9800 ;
      RECT 2.0400 0.6600 2.4500 0.7500 ;
      RECT 4.1050 0.6600 4.8150 0.7500 ;
      RECT 4.6800 1.2850 4.8400 1.7400 ;
      RECT 4.7300 0.9300 4.8400 1.2850 ;
      RECT 4.7300 0.8400 5.2800 0.9300 ;
      RECT 5.1750 0.9300 5.2800 0.9700 ;
      RECT 4.9250 0.6600 5.0950 0.8400 ;
      RECT 5.1750 0.9700 5.5200 1.0700 ;
      RECT 5.6400 1.0050 6.8850 1.1050 ;
      RECT 5.4100 1.2700 5.5100 1.5000 ;
      RECT 5.4100 1.1700 5.7400 1.2700 ;
      RECT 5.6400 1.1050 5.7400 1.1700 ;
      RECT 5.6400 0.8750 5.7400 1.0050 ;
      RECT 5.4100 0.7750 5.7400 0.8750 ;
      RECT 5.4100 0.6600 5.5100 0.7750 ;
      RECT 1.7050 0.4800 7.2950 0.5700 ;
      RECT 7.2050 0.5700 7.2950 0.9900 ;
      RECT 7.2050 0.9900 7.4950 1.0900 ;
      RECT 1.0650 0.8050 1.1650 1.2900 ;
      RECT 1.0650 1.2900 1.5250 1.3800 ;
      RECT 1.0650 0.7150 1.7950 0.8050 ;
      RECT 1.7050 0.5700 1.7950 0.7150 ;
      RECT 0.0500 1.8300 7.8700 1.9200 ;
      RECT 7.7800 1.1750 7.8700 1.8300 ;
      RECT 7.7800 0.9600 7.9150 1.1750 ;
      RECT 0.0500 1.5000 0.2050 1.8300 ;
      RECT 0.0500 0.9700 0.1400 1.5000 ;
      RECT 0.0500 0.6750 0.1400 0.8700 ;
      RECT 0.0500 0.5700 0.2100 0.6750 ;
      RECT 0.0500 0.8700 0.5550 0.9700 ;
      RECT 0.4550 0.9700 0.5550 1.0650 ;
      RECT 0.0500 0.4800 1.3000 0.5700 ;
      RECT 7.3900 0.5600 8.1000 0.6500 ;
      RECT 7.9250 0.5400 8.1000 0.5600 ;
      RECT 7.5850 0.7400 8.6000 0.8300 ;
      RECT 8.4250 0.6700 8.6000 0.7400 ;
      RECT 8.0050 1.4400 8.6100 1.5300 ;
      RECT 4.9600 1.6500 7.6750 1.7400 ;
      RECT 7.5850 0.8300 7.6750 1.6500 ;
      RECT 8.0050 0.8300 8.0950 1.4400 ;
      RECT 4.9600 1.0200 5.0600 1.6500 ;
      RECT 7.9650 1.6200 8.8900 1.7200 ;
      RECT 8.8000 1.1500 8.8900 1.6200 ;
      RECT 8.8000 1.0500 9.2250 1.1500 ;
      RECT 8.8000 0.5800 8.8900 1.0500 ;
      RECT 8.1900 0.4800 8.8900 0.5800 ;
      RECT 7.9650 1.7200 8.0750 1.9900 ;
      RECT 9.3150 1.0500 10.4850 1.1500 ;
      RECT 8.9950 1.4300 9.0950 1.9800 ;
      RECT 8.9950 0.4500 9.0950 0.8400 ;
      RECT 8.9950 1.3300 9.4150 1.4300 ;
      RECT 9.3150 1.1500 9.4150 1.3300 ;
      RECT 9.3150 0.9400 9.4150 1.0500 ;
      RECT 8.9950 0.8400 9.4150 0.9400 ;
  END
END BENC_X6M_A12TH

MACRO BENC_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 12.6450 2.7200 ;
        RECT 0.2800 2.0450 0.4900 2.0800 ;
        RECT 2.3350 2.0400 2.5550 2.0800 ;
        RECT 9.2750 1.8400 9.3850 2.0800 ;
        RECT 9.7900 1.8400 9.8900 2.0800 ;
        RECT 10.3400 1.7600 10.4400 2.0800 ;
        RECT 10.8600 1.7600 10.9600 2.0800 ;
        RECT 11.3800 1.7600 11.4800 2.0800 ;
        RECT 11.9000 1.7600 12.0000 2.0800 ;
        RECT 12.4200 1.7600 12.5200 2.0800 ;
    END
  END VDD

  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9850 1.5650 1.1900 ;
        RECT 1.4500 0.8950 2.0000 0.9850 ;
        RECT 1.9100 0.9850 2.0000 1.4700 ;
        RECT 1.9100 1.4700 4.8900 1.5600 ;
        RECT 4.7900 0.9550 4.8900 1.4700 ;
    END
    ANTENNAGATEAREA 0.2061 ;
  END M1

  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 1.1550 0.4300 1.3900 ;
        RECT 0.3300 1.3900 0.4300 1.6500 ;
        RECT 0.3300 1.6500 5.1050 1.7400 ;
        RECT 5.0050 1.1900 5.1050 1.6500 ;
        RECT 5.0050 0.9450 5.1500 1.1900 ;
    END
    ANTENNAGATEAREA 0.1617 ;
  END M0

  PIN X2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6550 0.8200 4.3650 0.9500 ;
        RECT 4.2350 0.9500 4.3650 1.2500 ;
        RECT 2.6550 0.7050 2.7550 0.8200 ;
        RECT 3.1750 0.7050 3.2750 0.8200 ;
        RECT 3.6950 0.7050 3.7950 0.8200 ;
        RECT 4.2150 0.7050 4.3150 0.8200 ;
        RECT 2.6200 1.2500 4.3650 1.3800 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END X2

  PIN AN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4150 1.2500 8.1850 1.4050 ;
        RECT 7.8350 0.9500 7.9650 1.2500 ;
        RECT 6.4700 0.8200 8.1300 0.9500 ;
        RECT 6.4700 0.7050 6.5700 0.8200 ;
        RECT 6.9900 0.7050 7.0900 0.8200 ;
        RECT 7.5100 0.7050 7.6100 0.8200 ;
        RECT 8.0300 0.7050 8.1300 0.8200 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END AN

  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.6000 1.2500 12.2600 1.3800 ;
        RECT 10.6000 1.3800 10.7000 1.7350 ;
        RECT 11.1200 1.3800 11.2200 1.7350 ;
        RECT 11.6400 1.3800 11.7400 1.7350 ;
        RECT 12.1600 1.3800 12.2600 1.7350 ;
        RECT 12.1300 0.9500 12.2600 1.2500 ;
        RECT 10.6000 0.8200 12.2600 0.9500 ;
        RECT 11.1200 0.4500 11.2200 0.8200 ;
        RECT 11.6400 0.4500 11.7400 0.8200 ;
        RECT 12.1600 0.4500 12.2600 0.8200 ;
        RECT 10.6000 0.4400 10.7000 0.8200 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END SN

  PIN M2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2500 1.0100 9.7500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0993 ;
  END M2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 12.6450 0.3200 ;
        RECT 4.8950 0.3200 5.1050 0.3750 ;
        RECT 8.7350 0.3200 8.8850 0.4550 ;
        RECT 10.3400 0.3200 10.4400 0.6400 ;
        RECT 10.8600 0.3200 10.9600 0.5750 ;
        RECT 11.3800 0.3200 11.4800 0.5750 ;
        RECT 11.9000 0.3200 12.0000 0.5750 ;
        RECT 12.4200 0.3200 12.5200 0.6400 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.5550 1.4400 0.7650 1.5600 ;
      RECT 0.6650 0.7750 0.7650 1.4400 ;
      RECT 0.5600 0.6600 0.7650 0.7750 ;
      RECT 0.8800 1.4700 1.8200 1.5600 ;
      RECT 1.7100 1.0750 1.8200 1.4700 ;
      RECT 0.8800 0.6800 0.9750 1.4700 ;
      RECT 2.3500 1.0500 3.8600 1.1500 ;
      RECT 2.0900 1.2700 2.4500 1.3800 ;
      RECT 2.3500 1.1500 2.4500 1.2700 ;
      RECT 2.3500 0.7500 2.4500 1.0500 ;
      RECT 2.0400 0.6600 2.4500 0.7500 ;
      RECT 4.6350 0.6600 5.3450 0.7500 ;
      RECT 5.2100 1.2850 5.3700 1.7400 ;
      RECT 5.2600 0.9300 5.3700 1.2850 ;
      RECT 5.2600 0.8400 5.8100 0.9300 ;
      RECT 5.7050 0.9300 5.8100 0.9700 ;
      RECT 5.4700 0.6800 5.5700 0.8400 ;
      RECT 5.7050 0.9700 6.0500 1.0700 ;
      RECT 6.1700 1.0500 7.6300 1.1500 ;
      RECT 5.9400 1.2700 6.0400 1.5000 ;
      RECT 5.9400 1.1700 6.2700 1.2700 ;
      RECT 6.1700 1.1500 6.2700 1.1700 ;
      RECT 6.1700 0.8750 6.2700 1.0500 ;
      RECT 5.9400 0.7750 6.2700 0.8750 ;
      RECT 5.9400 0.6600 6.0400 0.7750 ;
      RECT 1.7050 0.4800 8.3400 0.5700 ;
      RECT 8.2500 0.5700 8.3400 0.9900 ;
      RECT 8.2500 0.9900 8.5500 1.0900 ;
      RECT 1.0650 0.8050 1.1650 1.2900 ;
      RECT 1.0650 1.2900 1.5250 1.3800 ;
      RECT 1.0650 0.7150 1.7950 0.8050 ;
      RECT 1.7050 0.5700 1.7950 0.7150 ;
      RECT 0.0500 1.8300 8.7450 1.9200 ;
      RECT 8.6250 1.5600 8.7450 1.8300 ;
      RECT 8.6250 1.4600 8.9250 1.5600 ;
      RECT 8.8350 1.1750 8.9250 1.4600 ;
      RECT 8.8350 0.9650 8.9700 1.1750 ;
      RECT 0.0500 1.5000 0.2050 1.8300 ;
      RECT 0.0500 0.9700 0.1400 1.5000 ;
      RECT 0.0500 0.6750 0.1400 0.8700 ;
      RECT 0.0500 0.5700 0.2100 0.6750 ;
      RECT 0.0500 0.8700 0.5550 0.9700 ;
      RECT 0.4550 0.9700 0.5550 1.0650 ;
      RECT 0.0500 0.4800 1.2800 0.5700 ;
      RECT 8.4450 0.5600 9.1550 0.6500 ;
      RECT 8.9800 0.5400 9.1550 0.5600 ;
      RECT 8.6400 0.7400 9.6550 0.8300 ;
      RECT 9.4800 0.6700 9.6550 0.7400 ;
      RECT 9.0600 1.3000 9.4550 1.3900 ;
      RECT 9.3650 1.3900 9.4550 1.4550 ;
      RECT 9.3650 1.4550 9.6650 1.5450 ;
      RECT 5.4900 1.6500 8.4550 1.7400 ;
      RECT 8.3500 1.3500 8.4550 1.6500 ;
      RECT 8.3500 1.2500 8.7300 1.3500 ;
      RECT 8.6400 0.8300 8.7300 1.2500 ;
      RECT 9.0600 0.8300 9.1500 1.3000 ;
      RECT 5.4900 1.0200 5.5900 1.6500 ;
      RECT 8.9850 1.6500 9.9450 1.7500 ;
      RECT 9.8550 1.1500 9.9450 1.6500 ;
      RECT 9.8550 1.0500 10.2900 1.1500 ;
      RECT 9.8550 0.5800 9.9450 1.0500 ;
      RECT 9.2450 0.4800 9.9450 0.5800 ;
      RECT 8.9850 1.7500 9.1550 1.9900 ;
      RECT 10.4000 1.0500 11.8850 1.1500 ;
      RECT 10.0500 1.3500 10.1500 1.8800 ;
      RECT 10.0500 0.4500 10.1500 0.7700 ;
      RECT 10.0500 1.2500 10.5000 1.3500 ;
      RECT 10.4000 1.1500 10.5000 1.2500 ;
      RECT 10.4000 0.8700 10.5000 1.0500 ;
      RECT 10.0500 0.7700 10.5000 0.8700 ;
  END
END BENC_X8M_A12TH

MACRO BMXIT_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 3.9250 1.7450 4.0250 2.0800 ;
        RECT 0.0750 1.5000 0.1750 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0000 1.3500 1.1000 ;
        RECT 1.1950 1.1000 1.3500 1.2700 ;
        RECT 1.2500 1.2700 1.3500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0576 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9400 0.2750 1.1400 ;
        RECT 0.0500 1.1400 0.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END AN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9500 1.2050 ;
        RECT 2.6500 1.2050 2.9500 1.3700 ;
        RECT 2.6500 1.3700 2.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0576 ;
  END X2

  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.7100 4.3500 1.5500 ;
        RECT 4.1850 1.5500 4.3500 1.6650 ;
        RECT 4.1850 0.6100 4.3500 0.7100 ;
        RECT 4.1850 1.6650 4.2850 1.9900 ;
        RECT 4.1850 0.4900 4.2850 0.6100 ;
    END
    ANTENNADIFFAREA 0.1848 ;
  END PPN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0050 1.5500 1.4650 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END SN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8300 ;
        RECT 2.6200 0.3200 2.7900 0.6450 ;
        RECT 3.8700 0.3200 4.0800 0.3800 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8100 2.7500 0.9900 ;
    END
    ANTENNAGATEAREA 0.0576 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 1.0400 0.6950 1.2550 0.7950 ;
      RECT 0.9600 1.3850 1.1600 1.5600 ;
      RECT 0.9600 1.0250 1.0500 1.3850 ;
      RECT 0.9600 0.9350 1.1300 1.0250 ;
      RECT 1.0400 0.7950 1.1300 0.9350 ;
      RECT 0.7800 1.6500 1.7700 1.7400 ;
      RECT 1.5900 1.5500 1.7700 1.6500 ;
      RECT 1.6800 0.7500 1.7700 1.5500 ;
      RECT 1.5600 0.6600 1.7700 0.7500 ;
      RECT 0.7800 0.8450 0.8700 1.6500 ;
      RECT 0.7800 0.6600 0.9500 0.8450 ;
      RECT 0.3350 0.5400 2.1600 0.5700 ;
      RECT 2.0700 0.5700 2.1600 1.4400 ;
      RECT 0.3350 0.4800 2.2900 0.5400 ;
      RECT 2.0700 1.4400 2.2800 1.5500 ;
      RECT 2.0450 0.4300 2.2900 0.4800 ;
      RECT 0.3350 1.5750 0.4650 1.8200 ;
      RECT 0.3750 0.8300 0.4650 1.5750 ;
      RECT 0.3350 0.5700 0.4650 0.8300 ;
      RECT 2.3900 1.3500 2.4800 1.5300 ;
      RECT 2.2500 1.2600 2.4800 1.3500 ;
      RECT 2.2500 0.6300 2.4800 0.7200 ;
      RECT 2.3900 0.4750 2.4800 0.6300 ;
      RECT 2.2500 0.7200 2.3400 1.2600 ;
      RECT 2.8650 1.4600 3.1500 1.5500 ;
      RECT 3.0600 0.9000 3.1500 1.4600 ;
      RECT 2.9250 0.8000 3.1500 0.9000 ;
      RECT 2.9250 0.4750 3.0250 0.8000 ;
      RECT 1.8700 1.6400 3.3300 1.7400 ;
      RECT 3.2400 0.7100 3.3300 1.6400 ;
      RECT 3.1350 0.5700 3.3300 0.7100 ;
      RECT 1.8700 0.6600 1.9800 1.6400 ;
      RECT 0.6000 1.8300 3.7700 1.9200 ;
      RECT 3.6800 1.5250 3.7700 1.8300 ;
      RECT 3.6450 1.4350 3.7700 1.5250 ;
      RECT 3.6450 0.7700 3.7350 1.4350 ;
      RECT 3.6450 0.6600 3.8400 0.7700 ;
      RECT 0.6000 0.6800 0.6900 1.8300 ;
      RECT 3.4200 1.5050 3.5550 1.7200 ;
      RECT 3.4650 0.7650 3.5550 1.5050 ;
      RECT 3.4200 0.5700 3.5550 0.7650 ;
      RECT 3.4200 0.4800 4.0950 0.5700 ;
      RECT 4.0050 0.5700 4.0950 1.4500 ;
  END
END BMXIT_X0P7M_A12TH

MACRO BMXIT_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 3.9100 1.7450 4.0100 2.0800 ;
        RECT 0.0750 1.5350 0.1750 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0000 1.3500 1.1000 ;
        RECT 1.1950 1.1000 1.3500 1.2700 ;
        RECT 1.2500 1.2700 1.3500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0705 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9400 0.2750 1.1400 ;
        RECT 0.0500 1.1400 0.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END AN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9500 1.2050 ;
        RECT 2.6500 1.2050 2.9500 1.3700 ;
        RECT 2.6500 1.3700 2.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0705 ;
  END X2

  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.8550 4.3500 1.3000 ;
        RECT 4.1700 1.3000 4.3500 1.4000 ;
        RECT 4.1700 0.7550 4.3500 0.8550 ;
        RECT 4.1700 1.4000 4.2700 1.7900 ;
        RECT 4.1700 0.4400 4.2700 0.7550 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END PPN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0050 1.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END SN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7850 ;
        RECT 2.6200 0.3200 2.7900 0.6450 ;
        RECT 3.8750 0.3200 4.0450 0.3800 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8100 2.7500 0.9900 ;
    END
    ANTENNAGATEAREA 0.0705 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 1.0400 0.6950 1.2550 0.7950 ;
      RECT 0.9600 1.3850 1.1600 1.5600 ;
      RECT 0.9600 1.0250 1.0500 1.3850 ;
      RECT 0.9600 0.9350 1.1300 1.0250 ;
      RECT 1.0400 0.7950 1.1300 0.9350 ;
      RECT 0.7800 1.6500 1.7700 1.7400 ;
      RECT 1.5900 1.6100 1.7700 1.6500 ;
      RECT 1.6800 0.7500 1.7700 1.6100 ;
      RECT 1.5600 0.6600 1.7700 0.7500 ;
      RECT 0.7800 0.8450 0.8700 1.6500 ;
      RECT 0.7800 0.6600 0.9500 0.8450 ;
      RECT 0.3350 0.5400 2.1600 0.5700 ;
      RECT 2.0700 0.5700 2.1600 1.4400 ;
      RECT 0.3350 0.4800 2.2900 0.5400 ;
      RECT 2.0700 1.4400 2.2800 1.5500 ;
      RECT 2.0450 0.4300 2.2900 0.4800 ;
      RECT 0.3350 1.5750 0.4650 1.9900 ;
      RECT 0.3750 0.7850 0.4650 1.5750 ;
      RECT 0.3350 0.5700 0.4650 0.7850 ;
      RECT 2.3900 1.3500 2.4800 1.5300 ;
      RECT 2.2500 1.2600 2.4800 1.3500 ;
      RECT 2.2500 0.6300 2.4800 0.7200 ;
      RECT 2.3900 0.4750 2.4800 0.6300 ;
      RECT 2.2500 0.7200 2.3400 1.2600 ;
      RECT 2.8650 1.4600 3.1500 1.5500 ;
      RECT 3.0600 0.8850 3.1500 1.4600 ;
      RECT 2.9250 0.7850 3.1500 0.8850 ;
      RECT 2.9250 0.4750 3.0250 0.7850 ;
      RECT 1.8700 1.6400 3.3300 1.7400 ;
      RECT 3.2400 0.6850 3.3300 1.6400 ;
      RECT 3.1600 0.4750 3.3300 0.6850 ;
      RECT 1.8700 0.6600 1.9800 1.6400 ;
      RECT 0.6000 1.8300 3.7700 1.9200 ;
      RECT 3.6800 1.5250 3.7700 1.8300 ;
      RECT 3.6450 1.4350 3.7700 1.5250 ;
      RECT 3.6450 0.7800 3.7350 1.4350 ;
      RECT 3.6450 0.6700 3.8400 0.7800 ;
      RECT 0.6000 0.6800 0.6900 1.8300 ;
      RECT 3.4200 1.5050 3.5550 1.7150 ;
      RECT 3.4650 0.7650 3.5550 1.5050 ;
      RECT 3.4200 0.5800 3.5550 0.7650 ;
      RECT 3.4200 0.4900 4.0350 0.5800 ;
      RECT 3.9450 0.5800 4.0350 1.2350 ;
  END
END BMXIT_X1M_A12TH

MACRO BMXIT_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.0750 1.6400 0.1750 2.0800 ;
        RECT 3.9000 1.6050 4.0000 2.0800 ;
        RECT 4.4250 1.6050 4.5250 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0000 1.3500 1.1000 ;
        RECT 1.1950 1.1000 1.3500 1.2700 ;
        RECT 1.2500 1.2700 1.3500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0888 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9400 0.2750 1.1400 ;
        RECT 0.0500 1.1400 0.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END AN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9500 1.2100 ;
        RECT 2.6500 1.2100 2.9500 1.3700 ;
        RECT 2.6500 1.3700 2.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0888 ;
  END X2

  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9500 4.5500 1.2500 ;
        RECT 4.1600 1.2500 4.5500 1.3500 ;
        RECT 4.1600 0.8500 4.5500 0.9500 ;
        RECT 4.1600 1.3500 4.2600 1.8750 ;
        RECT 4.1600 0.4900 4.2600 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END PPN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0050 1.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0711 ;
  END SN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8500 ;
        RECT 4.4250 0.3200 4.5250 0.6550 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8100 2.7500 0.9900 ;
    END
    ANTENNAGATEAREA 0.0888 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 1.0400 0.6950 1.2550 0.7950 ;
      RECT 0.9600 1.3850 1.1600 1.5600 ;
      RECT 0.9600 1.0250 1.0500 1.3850 ;
      RECT 0.9600 0.9350 1.1300 1.0250 ;
      RECT 1.0400 0.7950 1.1300 0.9350 ;
      RECT 0.7800 1.6500 1.7700 1.7400 ;
      RECT 1.6800 0.7500 1.7700 1.6500 ;
      RECT 1.5600 0.6600 1.7700 0.7500 ;
      RECT 0.7800 0.8450 0.8700 1.6500 ;
      RECT 0.7800 0.6600 0.9500 0.8450 ;
      RECT 0.3350 0.5400 2.1600 0.5700 ;
      RECT 2.0700 0.5700 2.1600 1.4400 ;
      RECT 0.3350 0.4800 2.2900 0.5400 ;
      RECT 2.0700 1.4400 2.2800 1.5500 ;
      RECT 2.0450 0.4300 2.2900 0.4800 ;
      RECT 0.3350 1.5750 0.4650 1.9900 ;
      RECT 0.3750 0.8700 0.4650 1.5750 ;
      RECT 0.3350 0.5700 0.4650 0.8700 ;
      RECT 2.3800 1.3500 2.4700 1.5300 ;
      RECT 2.2500 1.2600 2.4700 1.3500 ;
      RECT 2.2500 0.6300 2.4700 0.7200 ;
      RECT 2.3800 0.4750 2.4700 0.6300 ;
      RECT 2.2500 0.7200 2.3400 1.2600 ;
      RECT 2.8550 1.4600 3.1400 1.5500 ;
      RECT 3.0500 0.8850 3.1400 1.4600 ;
      RECT 2.9150 0.7850 3.1400 0.8850 ;
      RECT 2.9150 0.4750 3.0150 0.7850 ;
      RECT 1.8700 1.6400 3.3200 1.7400 ;
      RECT 3.2300 0.6850 3.3200 1.6400 ;
      RECT 3.1500 0.4750 3.3200 0.6850 ;
      RECT 1.8700 0.6600 1.9800 1.6400 ;
      RECT 0.6000 1.8300 3.7600 1.9200 ;
      RECT 3.6700 1.5100 3.7600 1.8300 ;
      RECT 3.6350 1.4200 3.7600 1.5100 ;
      RECT 3.6350 0.7800 3.7250 1.4200 ;
      RECT 3.6350 0.6700 3.8300 0.7800 ;
      RECT 0.6000 0.6800 0.6900 1.8300 ;
      RECT 3.9350 1.0500 4.2750 1.1500 ;
      RECT 3.4100 0.4900 4.0250 0.5800 ;
      RECT 3.9350 0.5800 4.0250 1.0500 ;
      RECT 3.4100 1.4400 3.5450 1.6750 ;
      RECT 3.4550 0.7650 3.5450 1.4400 ;
      RECT 3.4100 0.5800 3.5450 0.7650 ;
  END
END BMXIT_X1P4M_A12TH

MACRO BMXIT_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 0.0700 1.7600 0.1800 2.0800 ;
        RECT 4.6250 1.7600 4.7250 2.0800 ;
    END
  END VDD

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1650 1.0500 1.3900 1.2400 ;
        RECT 1.2500 1.2400 1.3900 1.3900 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END D1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.5250 ;
        RECT 4.6250 0.3200 4.7250 0.6400 ;
    END
  END VSS

  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.9500 4.7500 1.2500 ;
        RECT 4.3650 1.2500 4.7500 1.3500 ;
        RECT 4.3650 0.8500 4.7500 0.9500 ;
        RECT 4.3650 1.3500 4.4650 1.7400 ;
        RECT 4.3650 0.4400 4.4650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END PPN

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 0.6500 1.6150 0.9600 ;
        RECT 1.5050 0.9600 1.6150 1.0400 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END AN

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4100 1.0450 2.7900 1.1600 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END D0

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0750 1.0300 3.5950 1.1500 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END X2

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8100 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0846 ;
  END SN
  OBS
    LAYER M1 ;
      RECT 0.9650 0.8600 1.2050 0.9500 ;
      RECT 1.0950 0.6600 1.2050 0.8600 ;
      RECT 1.0650 1.4200 1.1550 1.5600 ;
      RECT 0.8200 1.3300 1.1550 1.4200 ;
      RECT 0.8200 1.2400 1.0750 1.3300 ;
      RECT 0.9650 0.9500 1.0750 1.2400 ;
      RECT 1.9050 0.6600 2.5350 0.7500 ;
      RECT 2.2950 0.7500 2.5350 0.7700 ;
      RECT 0.3450 0.4800 1.9950 0.5600 ;
      RECT 1.6600 0.5600 1.9950 0.5700 ;
      RECT 1.3200 0.4700 1.7050 0.4800 ;
      RECT 1.9050 0.5700 1.9950 0.6600 ;
      RECT 1.9050 0.7500 1.9950 1.4300 ;
      RECT 1.8050 1.4300 1.9950 1.5400 ;
      RECT 0.3450 0.5600 1.3650 0.5700 ;
      RECT 0.2800 1.8700 0.4950 1.9600 ;
      RECT 0.2800 1.6700 0.3700 1.8700 ;
      RECT 0.0450 1.5800 0.3700 1.6700 ;
      RECT 0.0450 0.6250 0.4350 0.7150 ;
      RECT 0.3450 0.5700 0.4350 0.6250 ;
      RECT 0.0450 0.7150 0.1350 1.5800 ;
      RECT 0.8050 1.6500 2.5450 1.7400 ;
      RECT 1.6250 1.3150 1.7150 1.6500 ;
      RECT 1.6250 1.2250 1.8150 1.3150 ;
      RECT 1.7050 0.6600 1.8150 1.2250 ;
      RECT 0.8050 1.6000 0.8950 1.6500 ;
      RECT 0.6400 1.5100 0.8950 1.6000 ;
      RECT 0.6400 1.1500 0.7300 1.5100 ;
      RECT 0.6400 1.0600 0.8750 1.1500 ;
      RECT 0.7850 0.7700 0.8750 1.0600 ;
      RECT 0.7850 0.6600 0.9950 0.7700 ;
      RECT 2.5650 1.3400 2.7750 1.3800 ;
      RECT 2.2250 1.2500 2.7750 1.3400 ;
      RECT 2.2250 0.8600 2.7350 0.9500 ;
      RECT 2.6250 0.6600 2.7350 0.8600 ;
      RECT 2.2250 0.9500 2.3150 1.2500 ;
      RECT 2.0850 1.4700 3.5400 1.5600 ;
      RECT 2.0850 0.4800 3.4700 0.5700 ;
      RECT 3.3800 0.5700 3.4700 0.6900 ;
      RECT 2.8950 0.5700 2.9850 1.4700 ;
      RECT 2.0850 1.4500 2.2700 1.4700 ;
      RECT 2.0850 0.4600 2.3050 0.4800 ;
      RECT 3.0750 1.2900 3.9050 1.3800 ;
      RECT 3.0750 1.2700 3.2950 1.2900 ;
      RECT 3.8050 0.9400 3.9050 1.2900 ;
      RECT 3.6850 0.9100 3.9050 0.9400 ;
      RECT 3.1450 0.8400 3.9050 0.9100 ;
      RECT 3.1450 0.8200 3.7500 0.8400 ;
      RECT 3.1450 0.6600 3.2350 0.8200 ;
      RECT 0.6050 1.8300 3.4200 1.9200 ;
      RECT 3.3300 1.7400 3.4200 1.8300 ;
      RECT 3.3300 1.6500 4.0850 1.7400 ;
      RECT 3.9950 0.7500 4.0850 1.6500 ;
      RECT 3.8250 0.6600 4.0850 0.7500 ;
      RECT 0.6050 1.7800 0.6950 1.8300 ;
      RECT 0.4600 1.6900 0.6950 1.7800 ;
      RECT 0.4600 0.9700 0.5500 1.6900 ;
      RECT 0.4600 0.8800 0.6950 0.9700 ;
      RECT 0.5850 0.6800 0.6950 0.8800 ;
      RECT 4.1750 1.0500 4.5200 1.1500 ;
      RECT 3.5800 1.8300 4.2650 1.9200 ;
      RECT 4.1750 1.1500 4.2650 1.8300 ;
      RECT 4.1750 0.5700 4.2650 1.0500 ;
      RECT 3.5700 0.4800 4.2650 0.5700 ;
  END
END BMXIT_X2M_A12TH

MACRO BMXT_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 4.2550 2.0100 4.4600 2.0800 ;
        RECT 0.0750 1.6150 0.1750 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0000 1.3500 1.1000 ;
        RECT 1.1950 1.1000 1.3500 1.2700 ;
        RECT 1.2500 1.2700 1.3500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0525 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9400 0.2750 1.1400 ;
        RECT 0.0500 1.1400 0.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END AN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9550 1.2100 ;
        RECT 2.6500 1.2100 2.9550 1.3700 ;
        RECT 2.6500 1.3700 2.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.054 ;
  END X2

  PIN PP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.7100 4.7500 1.4900 ;
        RECT 4.5700 1.4900 4.7500 1.5900 ;
        RECT 4.5800 0.6100 4.7500 0.7100 ;
        RECT 4.5700 1.5900 4.6700 1.9650 ;
        RECT 4.5800 0.4500 4.6800 0.6100 ;
    END
    ANTENNADIFFAREA 0.1899 ;
  END PP

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9250 1.5500 1.4150 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END SN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8250 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8100 2.7600 0.9900 ;
    END
    ANTENNAGATEAREA 0.0525 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 1.0400 0.6850 1.2550 0.7850 ;
      RECT 0.9600 1.3850 1.1600 1.5600 ;
      RECT 0.9600 1.0250 1.0500 1.3850 ;
      RECT 0.9600 0.9350 1.1300 1.0250 ;
      RECT 1.0400 0.7850 1.1300 0.9350 ;
      RECT 0.7800 1.6500 1.7700 1.7400 ;
      RECT 1.5900 1.5000 1.7700 1.6500 ;
      RECT 1.6800 0.7500 1.7700 1.5000 ;
      RECT 1.5600 0.6600 1.7700 0.7500 ;
      RECT 0.7800 0.8450 0.8700 1.6500 ;
      RECT 0.7800 0.6600 0.9500 0.8450 ;
      RECT 0.3350 0.5400 2.1600 0.5700 ;
      RECT 2.0700 0.5700 2.1600 1.4400 ;
      RECT 0.3350 0.4800 2.2900 0.5400 ;
      RECT 2.0700 1.4400 2.2800 1.5500 ;
      RECT 2.0450 0.4300 2.2900 0.4800 ;
      RECT 0.3350 1.6150 0.4650 1.8300 ;
      RECT 0.3750 0.8250 0.4650 1.6150 ;
      RECT 0.3350 0.5700 0.4650 0.8250 ;
      RECT 2.3800 1.3500 2.4700 1.5300 ;
      RECT 2.2500 1.2600 2.4700 1.3500 ;
      RECT 2.2500 0.6300 2.4800 0.7200 ;
      RECT 2.3900 0.4750 2.4800 0.6300 ;
      RECT 2.2500 0.7200 2.3400 1.2600 ;
      RECT 1.8700 1.6500 3.3200 1.7400 ;
      RECT 3.2300 1.0250 3.3200 1.6500 ;
      RECT 1.8700 0.6600 1.9800 1.6500 ;
      RECT 3.4200 0.8600 3.5100 1.7200 ;
      RECT 3.4000 0.6700 3.5100 0.8600 ;
      RECT 2.8650 1.4600 3.1400 1.5500 ;
      RECT 3.0500 0.8850 3.1400 1.4600 ;
      RECT 2.9250 0.7850 3.1400 0.8850 ;
      RECT 2.9250 0.5700 3.0250 0.7850 ;
      RECT 2.9250 0.4800 3.6900 0.5700 ;
      RECT 3.6000 0.5700 3.6900 1.1600 ;
      RECT 4.0400 0.6700 4.1300 1.7200 ;
      RECT 0.6000 1.8300 4.3100 1.9200 ;
      RECT 4.2200 0.9100 4.3100 1.8300 ;
      RECT 0.6000 0.6800 0.6900 1.8300 ;
      RECT 4.4000 0.9950 4.5600 1.2100 ;
      RECT 4.4000 0.5800 4.4900 0.9950 ;
      RECT 3.7800 0.4900 4.4900 0.5800 ;
      RECT 3.7800 0.5800 3.8700 1.7200 ;
  END
END BMXT_X0P7M_A12TH

MACRO BMXT_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 4.2750 2.0450 4.4450 2.0800 ;
        RECT 0.0750 1.5000 0.1750 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0000 1.3500 1.1000 ;
        RECT 1.1950 1.1000 1.3500 1.2700 ;
        RECT 1.2500 1.2700 1.3500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9400 0.2750 1.1400 ;
        RECT 0.0500 1.1400 0.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END AN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9550 1.2100 ;
        RECT 2.6500 1.2100 2.9550 1.3700 ;
        RECT 2.6500 1.3700 2.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END X2

  PIN PP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.8900 4.7500 1.4950 ;
        RECT 4.5700 1.4950 4.7500 1.5950 ;
        RECT 4.5800 0.7900 4.7500 0.8900 ;
        RECT 4.5700 1.5950 4.6700 1.9650 ;
        RECT 4.5800 0.4500 4.6800 0.7900 ;
    END
    ANTENNADIFFAREA 0.26715 ;
  END PP

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0050 1.5500 1.4700 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7800 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8100 2.7600 0.9900 ;
    END
    ANTENNAGATEAREA 0.0636 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 1.0400 0.6850 1.2550 0.7850 ;
      RECT 0.9600 1.3850 1.1600 1.5600 ;
      RECT 0.9600 1.0250 1.0500 1.3850 ;
      RECT 0.9600 0.9350 1.1300 1.0250 ;
      RECT 1.0400 0.7850 1.1300 0.9350 ;
      RECT 0.7800 1.6500 1.7700 1.7400 ;
      RECT 1.5900 1.5700 1.7700 1.6500 ;
      RECT 1.6800 0.7500 1.7700 1.5700 ;
      RECT 1.5600 0.6600 1.7700 0.7500 ;
      RECT 0.7800 0.8450 0.8700 1.6500 ;
      RECT 0.7800 0.6600 0.9500 0.8450 ;
      RECT 0.3350 0.5400 2.1600 0.5700 ;
      RECT 2.0700 0.5700 2.1600 1.4400 ;
      RECT 0.3350 0.4800 2.2900 0.5400 ;
      RECT 2.0700 1.4400 2.2800 1.5500 ;
      RECT 2.0450 0.4300 2.2900 0.4800 ;
      RECT 0.3350 1.6150 0.4650 1.8300 ;
      RECT 0.3750 0.7850 0.4650 1.6150 ;
      RECT 0.3350 0.5700 0.4650 0.7850 ;
      RECT 2.3800 1.3500 2.4700 1.5300 ;
      RECT 2.2500 1.2600 2.4700 1.3500 ;
      RECT 2.2500 0.6300 2.4800 0.7200 ;
      RECT 2.3900 0.4750 2.4800 0.6300 ;
      RECT 2.2500 0.7200 2.3400 1.2600 ;
      RECT 1.8700 1.6500 3.3200 1.7400 ;
      RECT 3.2300 1.0100 3.3200 1.6500 ;
      RECT 1.8700 0.6600 1.9800 1.6500 ;
      RECT 3.4200 0.8350 3.5100 1.6200 ;
      RECT 3.4000 0.6700 3.5100 0.8350 ;
      RECT 2.8650 1.4600 3.1400 1.5500 ;
      RECT 3.0500 0.8850 3.1400 1.4600 ;
      RECT 2.9250 0.7850 3.1400 0.8850 ;
      RECT 2.9250 0.5700 3.0250 0.7850 ;
      RECT 2.9250 0.4800 3.6900 0.5700 ;
      RECT 3.6000 0.5700 3.6900 1.1600 ;
      RECT 4.0400 0.6700 4.1300 1.6200 ;
      RECT 0.6000 1.8300 4.3100 1.9200 ;
      RECT 4.2200 0.9600 4.3100 1.8300 ;
      RECT 0.6000 0.6800 0.6900 1.8300 ;
      RECT 4.4000 0.9950 4.5600 1.2100 ;
      RECT 4.4000 0.5800 4.4900 0.9950 ;
      RECT 3.7800 0.4900 4.4900 0.5800 ;
      RECT 3.7800 0.5800 3.8700 1.6200 ;
  END
END BMXT_X1M_A12TH

MACRO BMXT_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 4.2650 2.0100 4.4350 2.0800 ;
        RECT 4.8250 1.6050 4.9250 2.0800 ;
        RECT 0.0750 1.5350 0.1750 2.0800 ;
    END
  END VDD

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0000 1.3500 1.1000 ;
        RECT 1.1950 1.1000 1.3500 1.2700 ;
        RECT 1.2500 1.2700 1.3500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9400 0.2750 1.1400 ;
        RECT 0.0500 1.1400 0.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END AN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 1.0100 2.9500 1.2100 ;
        RECT 2.6500 1.2100 2.9500 1.3700 ;
        RECT 2.6500 1.3700 2.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END X2

  PIN PP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.9500 4.9500 1.2500 ;
        RECT 4.5600 1.2500 4.9500 1.3500 ;
        RECT 4.5700 0.8500 4.9500 0.9500 ;
        RECT 4.5600 1.3500 4.6600 1.9450 ;
        RECT 4.5700 0.4500 4.6800 0.8500 ;
    END
    ANTENNADIFFAREA 0.236775 ;
  END PP

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 1.0050 1.5500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END SN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8500 ;
        RECT 4.8250 0.3200 4.9250 0.6550 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.8100 2.7500 0.9900 ;
    END
    ANTENNAGATEAREA 0.0822 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 1.0400 0.6850 1.2550 0.7850 ;
      RECT 0.9600 1.3850 1.1600 1.5600 ;
      RECT 0.9600 1.0250 1.0500 1.3850 ;
      RECT 0.9600 0.9350 1.1300 1.0250 ;
      RECT 1.0400 0.7850 1.1300 0.9350 ;
      RECT 0.7800 1.6500 1.7700 1.7400 ;
      RECT 1.6800 0.7500 1.7700 1.6500 ;
      RECT 1.5600 0.6600 1.7700 0.7500 ;
      RECT 0.7800 0.8450 0.8700 1.6500 ;
      RECT 0.7800 0.6600 0.9500 0.8450 ;
      RECT 0.3350 0.5400 2.1600 0.5700 ;
      RECT 2.0700 0.5700 2.1600 1.4400 ;
      RECT 0.3350 0.4800 2.2900 0.5400 ;
      RECT 2.0700 1.4400 2.2800 1.5500 ;
      RECT 2.0450 0.4300 2.2900 0.4800 ;
      RECT 0.3350 1.5750 0.4650 1.9900 ;
      RECT 0.3750 0.8700 0.4650 1.5750 ;
      RECT 0.3350 0.5700 0.4650 0.8700 ;
      RECT 2.3800 1.3500 2.4700 1.5300 ;
      RECT 2.2500 1.2600 2.4700 1.3500 ;
      RECT 2.2500 0.6300 2.4700 0.7200 ;
      RECT 2.3800 0.4750 2.4700 0.6300 ;
      RECT 2.2500 0.7200 2.3400 1.2600 ;
      RECT 1.8700 1.6500 3.3100 1.7400 ;
      RECT 3.2200 1.0100 3.3100 1.6500 ;
      RECT 1.8700 0.6600 1.9800 1.6500 ;
      RECT 3.4100 0.8350 3.5000 1.6200 ;
      RECT 3.3900 0.6700 3.5000 0.8350 ;
      RECT 2.8550 1.4600 3.1300 1.5500 ;
      RECT 3.0400 0.8850 3.1300 1.4600 ;
      RECT 2.9150 0.7850 3.1300 0.8850 ;
      RECT 2.9150 0.5700 3.0150 0.7850 ;
      RECT 2.9150 0.4800 3.6800 0.5700 ;
      RECT 3.5900 0.5700 3.6800 1.1500 ;
      RECT 4.0300 0.6700 4.1200 1.6200 ;
      RECT 0.6000 1.8300 4.3000 1.9200 ;
      RECT 4.2100 0.8900 4.3000 1.8300 ;
      RECT 0.6000 0.6800 0.6900 1.8300 ;
      RECT 4.3900 1.0500 4.6750 1.1500 ;
      RECT 4.3900 0.5800 4.4800 1.0500 ;
      RECT 3.7700 0.4900 4.4800 0.5800 ;
      RECT 3.7700 0.5800 3.8600 1.6200 ;
  END
END BMXT_X1P4M_A12TH

MACRO BMXT_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 1.3250 2.0100 1.4950 2.0800 ;
        RECT 5.2250 1.7600 5.3250 2.0800 ;
        RECT 0.0700 1.6850 0.1800 2.0800 ;
    END
  END VDD

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2350 0.8100 0.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0801 ;
  END SN

  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2400 1.0200 3.8400 1.1500 ;
        RECT 3.2400 1.1500 3.3550 1.1900 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END X2

  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4100 1.0450 2.7900 1.1600 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END D0

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 0.6500 1.6150 0.9600 ;
        RECT 1.5050 0.9600 1.6150 1.0200 ;
    END
    ANTENNAGATEAREA 0.0801 ;
  END AN

  PIN PP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 0.9500 5.3500 1.2500 ;
        RECT 4.9650 1.2500 5.3500 1.3500 ;
        RECT 4.9650 0.8500 5.3500 0.9500 ;
        RECT 4.9650 1.3500 5.0650 1.7000 ;
        RECT 4.9650 0.4450 5.0650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END PP

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.5250 ;
        RECT 3.3000 0.3200 3.4700 0.4050 ;
        RECT 5.2250 0.3200 5.3250 0.6400 ;
    END
  END VSS

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1650 1.0500 1.3900 1.2400 ;
        RECT 1.2500 1.2400 1.3900 1.3900 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END D1
  OBS
    LAYER M1 ;
      RECT 0.9650 0.8600 1.2050 0.9500 ;
      RECT 1.0950 0.6600 1.2050 0.8600 ;
      RECT 1.0500 1.4200 1.1400 1.5600 ;
      RECT 0.8200 1.3300 1.1400 1.4200 ;
      RECT 0.8200 1.2400 1.0750 1.3300 ;
      RECT 0.9650 0.9500 1.0750 1.2400 ;
      RECT 1.9050 0.6600 2.5350 0.7700 ;
      RECT 0.3450 0.4800 1.9950 0.5600 ;
      RECT 1.6600 0.5600 1.9950 0.5700 ;
      RECT 1.3100 0.4700 1.7050 0.4800 ;
      RECT 1.9050 0.5700 1.9950 0.6600 ;
      RECT 1.9750 0.7700 2.0650 1.2900 ;
      RECT 1.8250 1.2900 2.0650 1.3800 ;
      RECT 0.3450 0.5600 1.3550 0.5700 ;
      RECT 0.2800 1.8700 0.4750 1.9600 ;
      RECT 0.2800 1.5250 0.3700 1.8700 ;
      RECT 0.0450 1.4350 0.3700 1.5250 ;
      RECT 0.0450 0.6250 0.4350 0.7150 ;
      RECT 0.3450 0.5700 0.4350 0.6250 ;
      RECT 0.0450 0.7150 0.1350 1.4350 ;
      RECT 1.6250 1.4700 2.5450 1.5600 ;
      RECT 0.8050 1.6500 1.7150 1.7400 ;
      RECT 1.6250 1.5600 1.7150 1.6500 ;
      RECT 1.6250 1.2000 1.7150 1.4700 ;
      RECT 1.6250 1.1100 1.8150 1.2000 ;
      RECT 1.7050 0.6600 1.8150 1.1100 ;
      RECT 0.8050 1.6000 0.8950 1.6500 ;
      RECT 0.6400 1.5100 0.8950 1.6000 ;
      RECT 0.6400 1.1500 0.7300 1.5100 ;
      RECT 0.6400 1.0600 0.8750 1.1500 ;
      RECT 0.7850 0.7700 0.8750 1.0600 ;
      RECT 0.7850 0.6600 0.9950 0.7700 ;
      RECT 2.2250 1.2900 2.7900 1.3800 ;
      RECT 2.2250 0.8600 2.7350 0.9500 ;
      RECT 2.6250 0.6600 2.7350 0.8600 ;
      RECT 2.2250 0.9500 2.3150 1.2900 ;
      RECT 2.0450 1.6500 3.5200 1.7400 ;
      RECT 3.4300 1.3500 3.5200 1.6500 ;
      RECT 3.4300 1.2400 3.6750 1.3500 ;
      RECT 2.8800 0.5700 2.9700 1.6500 ;
      RECT 2.0850 0.4800 2.9700 0.5700 ;
      RECT 2.0850 0.4600 2.3050 0.4800 ;
      RECT 3.0600 1.4300 3.2950 1.5400 ;
      RECT 3.0600 0.8400 4.1250 0.9300 ;
      RECT 3.9300 0.9300 4.1250 0.9400 ;
      RECT 4.0250 0.9400 4.1250 1.2850 ;
      RECT 3.8550 1.2850 4.1250 1.3750 ;
      RECT 3.0600 0.9300 3.1500 1.4300 ;
      RECT 3.0600 0.6800 3.2350 0.8400 ;
      RECT 3.6350 1.4700 4.3050 1.5600 ;
      RECT 4.2150 0.7500 4.3050 1.4700 ;
      RECT 3.5450 0.6600 4.3050 0.7500 ;
      RECT 4.3950 0.7500 4.5050 1.5250 ;
      RECT 4.3950 0.6600 4.5700 0.7500 ;
      RECT 0.6050 1.8300 3.8400 1.9200 ;
      RECT 3.7300 1.7400 3.8400 1.8300 ;
      RECT 3.7300 1.6500 4.6850 1.7400 ;
      RECT 4.5950 1.0050 4.6850 1.6500 ;
      RECT 0.6050 1.7800 0.6950 1.8300 ;
      RECT 0.4600 1.6900 0.6950 1.7800 ;
      RECT 0.4600 0.9700 0.5500 1.6900 ;
      RECT 0.4600 0.8800 0.6950 0.9700 ;
      RECT 0.5850 0.6800 0.6950 0.8800 ;
      RECT 4.7850 1.0500 5.1200 1.1500 ;
      RECT 3.9850 1.8300 4.8750 1.9200 ;
      RECT 4.7850 1.1500 4.8750 1.8300 ;
      RECT 4.7850 0.5700 4.8750 1.0500 ;
      RECT 3.8500 0.4800 4.8750 0.5700 ;
  END
END BMXT_X2M_A12TH

MACRO BUFH_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.8450 0.3200 ;
        RECT 0.3650 0.3200 0.4650 0.5000 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8100 0.3500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8300 0.7500 1.4600 ;
        RECT 0.6300 1.4600 0.7500 1.8900 ;
        RECT 0.6300 0.4400 0.7500 0.8300 ;
    END
    ANTENNADIFFAREA 0.1848 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.8450 2.7200 ;
        RECT 0.3650 1.7000 0.4650 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5000 0.5400 1.5900 ;
      RECT 0.4500 0.7000 0.5400 1.5000 ;
      RECT 0.0750 0.6100 0.5400 0.7000 ;
      RECT 0.0750 1.5900 0.1750 1.9050 ;
      RECT 0.0750 0.4900 0.1700 0.6100 ;
  END
END BUFH_X0P7M_A12TH

MACRO AOI222_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.2450 0.3200 ;
        RECT 0.6550 0.3200 0.7550 0.6300 ;
        RECT 1.6000 0.3200 1.7700 0.5050 ;
        RECT 2.5800 0.3200 2.7500 0.5050 ;
        RECT 3.4300 0.3200 3.5300 0.5600 ;
        RECT 4.5000 0.3200 4.6000 0.6300 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1750 1.0500 1.3500 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9950 1.0500 3.1950 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7850 0.8500 2.9050 0.9500 ;
        RECT 1.7850 0.9500 1.8850 1.2400 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8400 1.0400 4.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END C0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5600 0.8500 4.9900 0.9500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3500 1.2500 4.8600 1.3500 ;
        RECT 3.7200 1.3500 3.8200 1.7200 ;
        RECT 4.2400 1.3500 4.3400 1.7200 ;
        RECT 4.7600 1.3500 4.8600 1.7200 ;
        RECT 3.3500 0.7500 3.4500 1.2500 ;
        RECT 1.0800 0.6500 4.1150 0.7500 ;
        RECT 1.0800 0.4500 1.2500 0.6500 ;
        RECT 2.1200 0.4500 2.2900 0.6500 ;
        RECT 3.9450 0.4500 4.1150 0.6500 ;
    END
    ANTENNADIFFAREA 0.897 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.2450 2.7200 ;
        RECT 0.3350 1.7700 0.4350 2.0800 ;
        RECT 0.8550 1.7700 0.9550 2.0800 ;
        RECT 1.3750 1.7700 1.4750 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 0.8500 1.5800 0.9500 ;
        RECT 1.4800 0.9500 1.5800 1.2400 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A1
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5000 3.3500 1.5900 ;
      RECT 1.6350 1.5900 1.7350 1.9300 ;
      RECT 0.0750 1.5900 0.1750 1.9300 ;
      RECT 0.5950 1.5900 0.6950 1.9300 ;
      RECT 1.1150 1.5900 1.2150 1.9300 ;
      RECT 1.8450 1.8300 5.1200 1.9200 ;
      RECT 5.0200 1.4900 5.1200 1.8300 ;
      RECT 3.4650 1.5100 3.5550 1.8300 ;
      RECT 3.9800 1.4500 4.0800 1.8300 ;
      RECT 4.5000 1.4900 4.6000 1.8300 ;
  END
END AOI222_X3M_A12TH

MACRO AOI222_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7650 ;
        RECT 1.0950 0.3200 1.2650 0.5550 ;
        RECT 2.1350 0.3200 2.3050 0.5550 ;
        RECT 3.1750 0.3200 3.3450 0.5550 ;
        RECT 4.2150 0.3200 4.3850 0.5550 ;
        RECT 4.4950 0.3200 4.6650 0.5550 ;
        RECT 5.5350 0.3200 5.7050 0.5550 ;
        RECT 6.6100 0.3200 6.7100 0.7750 ;
    END
  END VSS

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8950 1.0500 6.3400 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7500 4.5550 1.3450 ;
        RECT 4.4500 1.3450 6.5050 1.4450 ;
        RECT 0.6100 0.6500 6.2250 0.7500 ;
        RECT 0.6100 0.5400 0.7100 0.6500 ;
        RECT 1.6500 0.5400 1.7500 0.6500 ;
        RECT 2.6900 0.5400 2.7900 0.6500 ;
        RECT 3.7300 0.5400 3.8300 0.6500 ;
        RECT 5.0150 0.4350 5.1850 0.6500 ;
        RECT 6.0550 0.4350 6.2250 0.6500 ;
    END
    ANTENNADIFFAREA 1.196 ;
  END Y

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4500 0.9500 6.5500 1.2400 ;
        RECT 4.6850 0.8500 6.5500 0.9500 ;
        RECT 4.6850 0.9500 4.7850 1.2400 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END C1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5600 0.8500 3.9600 0.9500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 0.8500 1.8800 0.9500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2700 1.0500 4.2500 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.0500 2.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.8450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 1.3900 1.7700 1.4900 2.0800 ;
        RECT 1.9100 1.7700 2.0100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1700 1.6900 2.2700 1.9100 ;
      RECT 2.1700 1.6000 4.4050 1.6900 ;
      RECT 2.1700 1.5700 2.2700 1.6000 ;
      RECT 2.6900 1.2800 2.7900 1.6000 ;
      RECT 3.2100 1.2800 3.3100 1.6000 ;
      RECT 3.7300 1.2800 3.8300 1.6000 ;
      RECT 0.0900 1.4800 2.2700 1.5700 ;
      RECT 0.0900 1.5700 0.1900 1.9100 ;
      RECT 0.6100 1.5700 0.7100 1.9100 ;
      RECT 1.1300 1.5700 1.2300 1.9100 ;
      RECT 1.6500 1.5700 1.7500 1.9100 ;
      RECT 2.3750 1.8300 4.6500 1.9200 ;
      RECT 4.5100 1.6400 4.6500 1.8300 ;
      RECT 4.5100 1.5500 6.7100 1.6400 ;
      RECT 5.0500 1.6400 5.1500 1.9800 ;
      RECT 5.5700 1.6400 5.6700 1.9800 ;
      RECT 6.0900 1.6400 6.1900 1.9800 ;
      RECT 6.6100 1.6400 6.7100 1.9800 ;
  END
END AOI222_X4M_A12TH

MACRO AOI22_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.5700 ;
        RECT 1.1550 0.3200 1.3250 0.4950 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.6850 0.3500 1.1050 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 0.8500 0.9050 0.9500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.2500 0.7050 1.3500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.8000 1.1500 1.2200 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6900 1.3500 1.3400 ;
        RECT 0.9300 1.3400 1.3500 1.4400 ;
        RECT 0.6500 0.5900 1.3500 0.6900 ;
        RECT 0.9300 1.4400 1.0300 1.7200 ;
        RECT 0.6500 0.4450 0.7500 0.5900 ;
    END
    ANTENNADIFFAREA 0.165 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3650 1.6550 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6450 1.8300 1.2850 1.9200 ;
      RECT 1.1950 1.5500 1.2850 1.8300 ;
      RECT 0.0950 1.4750 0.7350 1.5650 ;
      RECT 0.6450 1.5650 0.7350 1.8300 ;
      RECT 0.0950 1.5650 0.1850 1.9700 ;
  END
END AOI22_X0P5M_A12TH

MACRO AOI22_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7050 ;
        RECT 1.1950 0.3200 1.2850 0.5000 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 0.8500 0.9100 0.9500 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.2500 0.7100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0850 0.8100 0.3550 0.9200 ;
        RECT 0.2450 0.9200 0.3550 1.1450 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.3450 ;
        RECT 0.9300 1.3450 1.3500 1.4450 ;
        RECT 0.6500 0.6000 1.3500 0.7000 ;
        RECT 0.9300 1.4450 1.0300 1.7100 ;
        RECT 0.6500 0.4900 0.7500 0.6000 ;
    END
    ANTENNADIFFAREA 0.2343 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.8250 1.1500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3650 1.7200 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6450 1.8300 1.2850 1.9200 ;
      RECT 1.1950 1.5500 1.2850 1.8300 ;
      RECT 0.0950 1.5100 0.7350 1.6000 ;
      RECT 0.6450 1.6000 0.7350 1.8300 ;
      RECT 0.0950 1.6000 0.1850 1.9450 ;
  END
END AOI22_X0P7M_A12TH

MACRO AOI22_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.6400 ;
        RECT 1.1800 0.3200 1.2800 0.6400 ;
    END
  END VSS

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7350 0.1600 1.1600 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.6900 0.5600 1.1200 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8850 0.9500 1.3050 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 0.8950 1.3500 1.3600 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.4300 0.7500 1.3000 ;
        RECT 0.3800 1.3000 0.7500 1.4000 ;
        RECT 0.3800 1.4000 0.4800 1.7100 ;
    END
    ANTENNADIFFAREA 0.3118 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.9200 1.7700 1.0200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6450 1.5000 1.2750 1.5900 ;
      RECT 1.1850 1.5900 1.2750 1.9200 ;
      RECT 0.1250 1.8300 0.7350 1.9200 ;
      RECT 0.6450 1.5900 0.7350 1.8300 ;
      RECT 0.1250 1.4900 0.2150 1.8300 ;
  END
END AOI22_X1M_A12TH

MACRO AOI22_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7550 ;
        RECT 1.1550 0.3200 1.2450 0.5550 ;
        RECT 2.1950 0.3200 2.2850 0.5550 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7600 2.3500 1.5600 ;
        RECT 1.3550 1.5600 2.3500 1.6600 ;
        RECT 0.9550 0.6600 2.3500 0.7600 ;
        RECT 0.9550 0.5800 1.0450 0.6600 ;
        RECT 0.5650 0.4800 1.0450 0.5800 ;
    END
    ANTENNADIFFAREA 0.426 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 0.8500 2.1400 0.9500 ;
        RECT 1.3150 0.9500 1.4150 1.0850 ;
        RECT 2.0400 0.9500 2.1400 1.3100 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 1.2400 1.9100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3600 1.7000 0.4500 2.0800 ;
        RECT 0.8900 1.7000 0.9800 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8500 1.1500 0.9500 ;
        RECT 0.2500 0.9500 0.3500 1.1150 ;
        RECT 1.0500 0.9500 1.1500 1.2750 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.2400 0.9050 1.3500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 1.1550 1.8300 2.3250 1.9200 ;
      RECT 1.1550 1.5900 1.2450 1.8300 ;
      RECT 0.0900 1.5000 1.2450 1.5900 ;
      RECT 0.0900 1.5900 0.1800 1.9250 ;
      RECT 0.6250 1.5900 0.7150 1.9300 ;
  END
END AOI22_X1P4M_A12TH

MACRO AOI22_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6200 ;
        RECT 1.1500 0.3200 1.2500 0.5700 ;
        RECT 2.1950 0.3200 2.2850 0.5700 ;
    END
  END VSS

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2550 0.8500 2.1350 0.9500 ;
        RECT 1.2550 0.9500 1.3550 1.1300 ;
        RECT 2.0350 0.9500 2.1350 1.0900 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7600 2.3500 1.3000 ;
        RECT 1.9300 1.3000 2.3500 1.4000 ;
        RECT 0.9500 0.6600 2.3500 0.7600 ;
        RECT 1.9300 1.4000 2.0300 1.6000 ;
        RECT 0.9500 0.5800 1.0400 0.6600 ;
        RECT 1.4100 1.6000 2.0300 1.7000 ;
        RECT 0.5650 0.4800 1.0400 0.5800 ;
        RECT 1.4100 1.3000 1.5100 1.6000 ;
    END
    ANTENNADIFFAREA 0.6 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0500 0.8600 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4850 1.0500 1.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 0.8500 1.1000 0.9600 ;
        RECT 0.9900 0.9600 1.1000 1.1050 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3600 1.7700 0.4500 2.0800 ;
        RECT 0.8900 1.7700 0.9800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1550 1.8300 2.3250 1.9200 ;
      RECT 1.1550 1.5750 1.2450 1.8300 ;
      RECT 0.0950 1.4850 1.2450 1.5750 ;
      RECT 0.0950 1.5750 0.1850 1.9150 ;
      RECT 0.6250 1.5750 0.7150 1.9150 ;
  END
END AOI22_X2M_A12TH

MACRO AOI22_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 1.1350 0.3200 1.2250 0.3700 ;
        RECT 1.6550 0.3200 1.7450 0.5700 ;
        RECT 2.1750 0.3200 2.2650 0.3700 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6700 1.0450 3.1150 1.1550 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8100 1.0500 2.2750 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0400 1.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.7800 2.5500 1.2500 ;
        RECT 1.9100 1.2500 3.0500 1.3500 ;
        RECT 0.0900 0.6800 3.3100 0.7800 ;
        RECT 1.9100 1.3500 2.0100 1.7200 ;
        RECT 2.4300 1.3500 2.5300 1.7200 ;
        RECT 2.9500 1.3500 3.0500 1.7200 ;
        RECT 0.0900 0.4100 0.1900 0.6800 ;
        RECT 3.2100 0.4100 3.3100 0.6800 ;
    END
    ANTENNADIFFAREA 0.9885 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0450 0.7200 1.1550 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.3100 0.4800 1.5450 0.5700 ;
      RECT 1.8550 0.4800 3.1000 0.5700 ;
      RECT 1.6550 1.8300 3.3050 1.9200 ;
      RECT 3.2150 1.4900 3.3050 1.8300 ;
      RECT 0.0950 1.4900 1.7450 1.5800 ;
      RECT 1.6550 1.5800 1.7450 1.8300 ;
      RECT 0.0950 1.5800 0.1850 1.9200 ;
      RECT 0.6150 1.5800 0.7050 1.9200 ;
      RECT 1.1350 1.5800 1.2250 1.9200 ;
      RECT 2.1750 1.5000 2.2650 1.8300 ;
      RECT 2.6950 1.5000 2.7850 1.8300 ;
  END
END AOI22_X3M_A12TH

MACRO AOI22_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.1350 0.3200 0.2250 0.6000 ;
        RECT 1.1750 0.3200 1.2650 0.5600 ;
        RECT 2.2150 0.3200 2.3050 0.5600 ;
        RECT 3.2650 0.3200 3.3550 0.5600 ;
        RECT 4.3050 0.3200 4.3950 0.6000 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 0.8500 1.9000 0.9350 ;
        RECT 0.5200 0.9350 1.9000 0.9500 ;
        RECT 0.5200 0.9500 0.8900 1.0350 ;
        RECT 1.5000 0.9500 1.9000 1.0050 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8900 0.8500 3.9900 0.9350 ;
        RECT 2.6100 0.9350 3.9900 0.9500 ;
        RECT 2.6100 0.9500 2.9800 1.0350 ;
        RECT 3.5950 0.9500 3.9900 1.0050 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 2.1300 1.3500 ;
        RECT 1.0400 1.0950 1.4100 1.2500 ;
        RECT 2.0400 1.0000 2.1300 1.2500 ;
        RECT 0.2400 0.9800 0.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2400 0.8000 4.3500 1.1250 ;
        RECT 2.4000 1.1250 4.3500 1.2150 ;
        RECT 3.1200 1.0950 3.4900 1.1250 ;
        RECT 2.4000 1.0000 2.4900 1.1250 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.6500 3.9150 0.7500 ;
        RECT 2.2200 0.7500 2.3100 1.3500 ;
        RECT 0.6150 0.4600 0.7850 0.6500 ;
        RECT 1.6550 0.4600 1.8250 0.6500 ;
        RECT 2.7050 0.4600 2.8750 0.6500 ;
        RECT 3.7450 0.4600 3.9150 0.6500 ;
        RECT 2.2200 1.3500 2.5750 1.4400 ;
        RECT 2.4850 1.4400 4.1350 1.5300 ;
        RECT 2.4850 1.5300 2.5750 1.7400 ;
        RECT 3.0050 1.5300 3.0950 1.7400 ;
        RECT 3.5250 1.5300 3.6150 1.7400 ;
        RECT 4.0450 1.5300 4.1350 1.7400 ;
        RECT 3.0050 1.3700 3.0950 1.4400 ;
        RECT 3.5250 1.3700 3.6150 1.4400 ;
        RECT 4.0450 1.3700 4.1350 1.4400 ;
    END
    ANTENNADIFFAREA 1.2 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 0.3950 1.7700 0.4850 2.0800 ;
        RECT 0.9150 1.7700 1.0050 2.0800 ;
        RECT 1.4350 1.7700 1.5250 2.0800 ;
        RECT 1.9550 1.7700 2.0450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2150 1.8300 4.3950 1.9200 ;
      RECT 4.3050 1.5500 4.3950 1.8300 ;
      RECT 2.2150 1.6300 2.3050 1.8300 ;
      RECT 0.1350 1.5300 2.3050 1.6300 ;
      RECT 2.7450 1.9200 2.8350 1.9900 ;
      RECT 2.7450 1.6200 2.8350 1.8300 ;
      RECT 3.2650 1.9200 3.3550 1.9900 ;
      RECT 3.2650 1.6200 3.3550 1.8300 ;
      RECT 3.7850 1.9200 3.8750 1.9900 ;
      RECT 3.7850 1.6200 3.8750 1.8300 ;
      RECT 0.1350 1.6300 0.2250 1.9600 ;
      RECT 0.6550 1.6300 0.7450 1.9600 ;
      RECT 1.1750 1.6300 1.2650 1.9600 ;
      RECT 1.6950 1.6300 1.7850 1.9600 ;
  END
END AOI22_X4M_A12TH

MACRO AOI22_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.1600 0.3200 0.2500 0.5600 ;
        RECT 0.7150 0.3200 0.8850 0.3950 ;
        RECT 1.3850 0.3200 1.5550 0.3950 ;
        RECT 5.1150 0.3200 5.2850 0.3900 ;
        RECT 5.6850 0.3200 5.8550 0.3900 ;
        RECT 6.2700 0.3200 6.3600 0.6150 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 1.0500 1.5150 1.1500 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0500 3.0650 1.1600 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7000 1.0500 4.5000 1.1600 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3000 1.0500 6.1000 1.1600 ;
    END
    ANTENNAGATEAREA 0.5406 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.2500 6.3000 1.3500 ;
        RECT 3.5300 1.3500 3.7000 1.5950 ;
        RECT 4.0500 1.3500 4.2200 1.5950 ;
        RECT 4.5700 1.3500 4.7400 1.5950 ;
        RECT 5.0900 1.3500 5.2600 1.6000 ;
        RECT 5.6100 1.3500 5.7800 1.6000 ;
        RECT 6.1300 1.3500 6.3000 1.6000 ;
        RECT 3.2500 0.9600 3.3500 1.2500 ;
        RECT 2.2300 0.8700 4.7400 0.9600 ;
        RECT 2.2300 0.6650 2.4000 0.8700 ;
        RECT 2.7500 0.6650 2.9200 0.8700 ;
        RECT 4.0500 0.6600 4.2200 0.8700 ;
        RECT 4.5700 0.6600 4.7400 0.8700 ;
        RECT 3.3100 0.5900 3.4000 0.8700 ;
    END
    ANTENNADIFFAREA 1.802 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.3000 1.8800 0.4700 2.0800 ;
        RECT 0.8200 1.8800 0.9900 2.0800 ;
        RECT 1.4050 1.8800 1.5750 2.0800 ;
        RECT 1.9700 1.8800 2.1400 2.0800 ;
        RECT 2.4900 1.8800 2.6600 2.0800 ;
        RECT 3.0100 1.8800 3.1800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4200 0.4850 3.1400 0.5750 ;
      RECT 3.0500 0.5750 3.1400 0.7800 ;
      RECT 3.0500 0.4100 3.1400 0.4850 ;
      RECT 0.4200 0.5750 0.5100 0.8000 ;
      RECT 1.0900 0.5750 1.1800 0.8000 ;
      RECT 1.7600 0.5750 1.8500 0.8000 ;
      RECT 2.0100 0.5750 2.1000 0.8550 ;
      RECT 0.4200 0.4300 0.5100 0.4850 ;
      RECT 1.0900 0.4300 1.1800 0.4850 ;
      RECT 1.7600 0.4300 1.8500 0.4850 ;
      RECT 2.5300 0.5750 2.6200 0.7800 ;
      RECT 2.5300 0.4100 2.6200 0.4850 ;
      RECT 3.5700 0.4800 6.1000 0.5700 ;
      RECT 4.8700 0.5700 4.9600 0.8500 ;
      RECT 5.4400 0.5700 5.5300 0.8500 ;
      RECT 6.0100 0.5700 6.1000 0.8500 ;
      RECT 3.5700 0.5700 3.6600 0.7800 ;
      RECT 3.8300 0.5700 3.9200 0.7800 ;
      RECT 3.5700 0.4100 3.6600 0.4800 ;
      RECT 3.8300 0.4100 3.9200 0.4800 ;
      RECT 4.3500 0.5700 4.4400 0.7800 ;
      RECT 4.3500 0.4100 4.4400 0.4800 ;
      RECT 0.0800 1.7000 6.5200 1.7900 ;
      RECT 6.4300 1.7900 6.5200 1.8700 ;
      RECT 6.4300 1.5000 6.5200 1.7000 ;
      RECT 0.0800 1.7900 0.1700 1.8700 ;
      RECT 0.6000 1.7900 0.6900 1.8700 ;
      RECT 1.1200 1.7900 1.2100 1.8700 ;
      RECT 1.7500 1.7900 1.8400 1.8700 ;
      RECT 2.2700 1.7900 2.3600 1.8700 ;
      RECT 2.7900 1.7900 2.8800 1.8700 ;
      RECT 3.3100 1.7900 3.4000 1.8700 ;
      RECT 0.0800 1.5000 0.1700 1.7000 ;
      RECT 0.6000 1.5000 0.6900 1.7000 ;
      RECT 1.1200 1.5000 1.2100 1.7000 ;
      RECT 1.7500 1.5000 1.8400 1.7000 ;
      RECT 2.2700 1.5000 2.3600 1.7000 ;
      RECT 2.7900 1.5000 2.8800 1.7000 ;
      RECT 3.3100 1.5000 3.4000 1.7000 ;
      RECT 3.8300 1.7900 3.9200 1.8700 ;
      RECT 3.8300 1.5000 3.9200 1.7000 ;
      RECT 4.3500 1.7900 4.4400 1.8700 ;
      RECT 4.3500 1.5000 4.4400 1.7000 ;
      RECT 4.8700 1.7900 4.9600 1.8700 ;
      RECT 4.8700 1.5000 4.9600 1.7000 ;
      RECT 5.3900 1.7900 5.4800 1.8700 ;
      RECT 5.3900 1.5000 5.4800 1.7000 ;
      RECT 5.9100 1.7900 6.0000 1.8700 ;
      RECT 5.9100 1.5000 6.0000 1.7000 ;
  END
END AOI22_X6M_A12TH

MACRO AOI22_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 8.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.5600 ;
        RECT 0.6200 0.3200 0.7900 0.3950 ;
        RECT 1.2600 0.3200 1.4300 0.3950 ;
        RECT 1.9000 0.3200 2.0700 0.3950 ;
        RECT 6.6450 0.3200 6.8150 0.3900 ;
        RECT 7.2150 0.3200 7.3850 0.3900 ;
        RECT 7.7850 0.3200 7.9550 0.3900 ;
        RECT 8.3700 0.3200 8.4600 0.7000 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 1.0500 1.7950 1.1500 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3000 1.0450 2.7250 1.1950 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1750 1.0800 6.1550 1.1800 ;
        RECT 5.4100 1.0500 5.5900 1.0800 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6850 1.0650 8.1850 1.1650 ;
        RECT 7.0100 1.0500 7.1900 1.0650 ;
    END
    ANTENNAGATEAREA 0.7203 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4900 1.4500 8.3000 1.5500 ;
        RECT 4.4900 1.5500 4.6600 1.6100 ;
        RECT 5.0100 1.5500 5.1800 1.6100 ;
        RECT 5.5300 1.5500 5.7000 1.6100 ;
        RECT 6.0500 1.5500 6.2200 1.6100 ;
        RECT 6.5700 1.5500 6.7400 1.6100 ;
        RECT 7.0900 1.5500 7.2600 1.6100 ;
        RECT 7.6100 1.5500 7.7800 1.6100 ;
        RECT 8.1300 1.5500 8.3000 1.6100 ;
        RECT 4.4900 1.3200 4.6600 1.4500 ;
        RECT 5.0100 1.3200 5.1800 1.4500 ;
        RECT 5.5300 1.3200 5.7000 1.4500 ;
        RECT 6.0500 1.3200 6.3350 1.4500 ;
        RECT 6.5700 1.3200 6.7400 1.4500 ;
        RECT 7.0900 1.3200 7.2600 1.4500 ;
        RECT 7.6100 1.3200 7.7800 1.4500 ;
        RECT 8.1300 1.3200 8.3000 1.4500 ;
        RECT 4.5700 1.0450 4.6600 1.3200 ;
        RECT 6.2450 0.9600 6.3350 1.3200 ;
        RECT 2.8150 0.9550 4.6600 1.0450 ;
        RECT 5.0600 0.8700 6.3350 0.9600 ;
        RECT 2.7300 0.6650 2.9050 0.9550 ;
        RECT 3.2500 0.6650 3.4200 0.9550 ;
        RECT 3.7700 0.6650 3.9400 0.9550 ;
        RECT 4.3300 0.6250 4.4200 0.9550 ;
        RECT 5.0600 0.6600 5.2300 0.8700 ;
        RECT 5.5800 0.6600 5.7500 0.8700 ;
        RECT 6.1000 0.6600 6.2700 0.8700 ;
    END
    ANTENNADIFFAREA 2.401 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 8.6450 2.7200 ;
        RECT 0.3000 1.8800 0.4700 2.0800 ;
        RECT 0.8200 1.8800 0.9900 2.0800 ;
        RECT 1.3400 1.8800 1.5100 2.0800 ;
        RECT 1.8700 1.8800 2.0400 2.0800 ;
        RECT 2.4100 1.8800 2.5800 2.0800 ;
        RECT 2.9300 1.8800 3.1000 2.0800 ;
        RECT 3.4500 1.8800 3.6200 2.0800 ;
        RECT 3.9700 1.8800 4.1400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 0.4850 4.1600 0.5750 ;
      RECT 4.0700 0.5750 4.1600 0.8550 ;
      RECT 0.3400 0.5750 0.4300 0.8950 ;
      RECT 0.9800 0.5750 1.0700 0.9000 ;
      RECT 1.6200 0.5750 1.7100 0.9000 ;
      RECT 2.2600 0.5750 2.3500 0.9000 ;
      RECT 2.5100 0.5750 2.6000 0.9000 ;
      RECT 3.0300 0.5750 3.1200 0.8550 ;
      RECT 3.5500 0.5750 3.6400 0.8550 ;
      RECT 4.5900 0.4800 8.2000 0.5700 ;
      RECT 6.4000 0.5700 6.4900 0.7800 ;
      RECT 6.9700 0.5700 7.0600 0.8900 ;
      RECT 7.5400 0.5700 7.6300 0.8900 ;
      RECT 8.1100 0.5700 8.2000 0.8900 ;
      RECT 6.4000 0.4100 6.4900 0.4800 ;
      RECT 4.5900 0.5700 4.6800 0.8500 ;
      RECT 4.8400 0.5700 4.9300 0.8900 ;
      RECT 5.3600 0.5700 5.4500 0.7800 ;
      RECT 5.3600 0.4100 5.4500 0.4800 ;
      RECT 5.8800 0.5700 5.9700 0.7800 ;
      RECT 5.8800 0.4100 5.9700 0.4800 ;
      RECT 0.0800 1.7000 8.5200 1.7900 ;
      RECT 8.4300 1.7900 8.5200 1.8700 ;
      RECT 8.4300 1.5000 8.5200 1.7000 ;
      RECT 4.2700 1.7900 4.3600 1.8700 ;
      RECT 4.2700 1.5000 4.3600 1.7000 ;
      RECT 4.7500 1.7900 4.9200 1.9300 ;
      RECT 4.7500 1.6400 4.9200 1.7000 ;
      RECT 5.2700 1.7900 5.4400 1.9300 ;
      RECT 5.2700 1.6400 5.4400 1.7000 ;
      RECT 5.7900 1.7900 5.9600 1.9300 ;
      RECT 5.7900 1.6400 5.9600 1.7000 ;
      RECT 6.3100 1.7900 6.4800 1.9300 ;
      RECT 6.3100 1.6400 6.4800 1.7000 ;
      RECT 6.8300 1.7900 7.0000 1.9300 ;
      RECT 6.8300 1.6400 7.0000 1.7000 ;
      RECT 7.3500 1.7900 7.5200 1.9300 ;
      RECT 7.3500 1.6400 7.5200 1.7000 ;
      RECT 7.8700 1.7900 8.0400 1.9300 ;
      RECT 7.8700 1.6400 8.0400 1.7000 ;
      RECT 0.0800 1.7900 0.1700 1.8700 ;
      RECT 0.0800 1.5000 0.1700 1.7000 ;
      RECT 0.6000 1.7900 0.6900 1.8700 ;
      RECT 0.6000 1.5000 0.6900 1.7000 ;
      RECT 1.1200 1.7900 1.2100 1.8700 ;
      RECT 1.1200 1.5000 1.2100 1.7000 ;
      RECT 1.6400 1.7900 1.7300 1.8700 ;
      RECT 1.6400 1.5000 1.7300 1.7000 ;
      RECT 2.1900 1.7900 2.2800 1.8700 ;
      RECT 2.1900 1.5000 2.2800 1.7000 ;
      RECT 2.7100 1.7900 2.8000 1.8700 ;
      RECT 2.7100 1.5000 2.8000 1.7000 ;
      RECT 3.2300 1.7900 3.3200 1.8700 ;
      RECT 3.2300 1.5000 3.3200 1.7000 ;
      RECT 3.7500 1.7900 3.8400 1.8700 ;
      RECT 3.7500 1.5000 3.8400 1.7000 ;
  END
END AOI22_X8M_A12TH

MACRO AOI2XB1_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1050 0.3200 0.1950 0.8850 ;
        RECT 0.3750 0.3200 0.4650 0.4800 ;
        RECT 1.2300 0.3200 1.3200 0.5600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7500 1.3500 1.6200 ;
        RECT 1.2300 1.6200 1.3500 1.7100 ;
        RECT 0.8950 0.6500 1.3500 0.7500 ;
        RECT 1.2300 1.7100 1.3200 1.9900 ;
        RECT 0.8950 0.4200 0.9850 0.6500 ;
    END
    ANTENNADIFFAREA 0.142925 ;
  END Y

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 1.0000 0.3500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.6100 0.7500 0.9000 ;
        RECT 0.6500 0.9000 0.9250 0.9900 ;
        RECT 0.8350 0.9900 0.9250 1.0950 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9800 1.1550 1.3900 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.7100 1.7250 0.8000 2.0800 ;
        RECT 0.1800 1.3050 0.2700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4600 1.0850 0.6950 1.2750 ;
      RECT 0.4400 1.2850 0.5500 1.4550 ;
      RECT 0.4600 1.2750 0.5500 1.2850 ;
      RECT 0.4600 0.8950 0.5500 1.0850 ;
      RECT 0.3650 0.8050 0.5500 0.8950 ;
      RECT 0.3650 0.6850 0.4550 0.8050 ;
      RECT 0.4500 1.5450 1.0600 1.6350 ;
      RECT 0.9700 1.6350 1.0600 1.9750 ;
      RECT 0.4500 1.6350 0.5400 1.9900 ;
  END
END AOI2XB1_X0P5M_A12TH

MACRO AOI2XB1_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6700 ;
        RECT 0.6300 0.3200 0.7300 0.4750 ;
        RECT 1.4200 0.3200 1.5200 0.4500 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8950 1.3500 1.3200 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END B0

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.8150 0.3550 1.2150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END A1N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8900 1.7950 0.9900 2.0800 ;
        RECT 0.0900 1.3700 0.1900 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.1500 1.1500 1.3900 ;
        RECT 0.9400 1.0500 1.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.7500 1.5500 1.5700 ;
        RECT 1.3700 1.5700 1.5500 1.9600 ;
        RECT 1.1000 0.6500 1.5500 0.7500 ;
        RECT 1.1000 0.4450 1.2000 0.6500 ;
    END
    ANTENNADIFFAREA 0.200125 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.3500 1.3300 0.8200 1.4300 ;
      RECT 0.7200 0.7200 0.8200 1.3300 ;
      RECT 0.3500 0.6200 0.8200 0.7200 ;
      RECT 0.3500 1.4300 0.4500 1.5800 ;
      RECT 0.3500 0.4550 0.4500 0.6200 ;
      RECT 0.6300 1.5500 1.2500 1.6400 ;
      RECT 1.1500 1.6400 1.2500 1.9800 ;
      RECT 0.6300 1.6400 0.7300 1.9800 ;
  END
END AOI2XB1_X0P7M_A12TH

MACRO AOI2XB1_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7000 ;
        RECT 0.5950 0.3200 0.7650 0.5300 ;
        RECT 1.4100 0.3200 1.5100 0.4400 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 0.9800 1.3500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END B0

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8200 0.3500 1.2250 ;
    END
    ANTENNAGATEAREA 0.0273 ;
  END A1N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.8900 1.7700 0.9900 2.0800 ;
        RECT 0.0900 1.3700 0.1900 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1100 0.9550 1.3900 ;
        RECT 0.8500 1.0100 1.1400 1.1100 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3850 1.5100 1.5500 1.9200 ;
        RECT 1.4500 0.7500 1.5500 1.5100 ;
        RECT 1.0550 0.6500 1.5500 0.7500 ;
        RECT 1.0550 0.4600 1.2250 0.6500 ;
    END
    ANTENNADIFFAREA 0.294375 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.3500 1.3450 0.7300 1.4350 ;
      RECT 0.6400 0.7200 0.7300 1.3450 ;
      RECT 0.3550 0.6300 0.7300 0.7200 ;
      RECT 0.3500 1.4350 0.4500 1.5550 ;
      RECT 0.3550 0.4650 0.4450 0.6300 ;
      RECT 0.6350 1.5500 1.2500 1.6400 ;
      RECT 1.1500 1.6400 1.2500 1.9800 ;
      RECT 0.6350 1.6400 0.7250 1.9800 ;
  END
END AOI2XB1_X1M_A12TH

MACRO AOI2XB1_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0850 0.3200 0.1950 0.6850 ;
        RECT 0.6400 0.3200 0.7500 0.7600 ;
        RECT 1.6800 0.3200 1.7900 0.5450 ;
        RECT 2.2150 0.3200 2.3250 0.5750 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.8100 0.3500 1.2400 ;
    END
    ANTENNAGATEAREA 0.0375 ;
  END A1N

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2400 0.7700 2.3500 1.1900 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9750 1.0500 1.4150 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 1.0900 2.0600 1.1900 ;
        RECT 1.9600 1.1900 2.0600 1.7150 ;
        RECT 1.8500 0.7500 1.9500 1.0900 ;
        RECT 1.1300 0.6500 2.0600 0.7500 ;
        RECT 1.1300 0.4600 1.3000 0.6500 ;
        RECT 1.9600 0.4200 2.0600 0.6500 ;
    END
    ANTENNADIFFAREA 0.266 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.9050 1.5150 1.0050 2.0800 ;
        RECT 1.4250 1.5150 1.5250 2.0800 ;
        RECT 0.0950 1.3400 0.1950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.7650 0.8600 1.6250 0.9500 ;
      RECT 1.5350 0.9500 1.6250 1.1900 ;
      RECT 0.4550 1.0500 0.8550 1.1500 ;
      RECT 0.7650 0.9500 0.8550 1.0500 ;
      RECT 0.3500 1.4850 0.4500 1.7850 ;
      RECT 0.3500 1.3850 0.5450 1.4850 ;
      RECT 0.4550 1.1500 0.5450 1.3850 ;
      RECT 0.4550 0.6600 0.5450 1.0500 ;
      RECT 0.3000 0.5600 0.5450 0.6600 ;
      RECT 1.6850 1.8200 2.3200 1.9200 ;
      RECT 2.2200 1.4850 2.3200 1.8200 ;
      RECT 1.6850 1.3900 1.7850 1.8200 ;
      RECT 0.6450 1.3000 1.7850 1.3900 ;
      RECT 0.6450 1.3900 0.7450 1.7300 ;
      RECT 1.1650 1.3900 1.2650 1.7300 ;
  END
END AOI2XB1_X1P4M_A12TH

MACRO AOI2XB1_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.8700 ;
        RECT 0.6350 0.3200 0.7450 0.6500 ;
        RECT 1.6450 0.3200 1.8150 0.5600 ;
        RECT 2.2150 0.3200 2.3150 0.6250 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9900 0.1600 1.4100 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9850 1.0500 1.4200 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.9000 1.7700 1.0000 2.0800 ;
        RECT 1.4200 1.7700 1.5200 2.0800 ;
        RECT 0.0900 1.5700 0.1900 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1250 0.6500 2.0500 0.7500 ;
        RECT 1.8550 0.7500 1.9450 1.2550 ;
        RECT 1.1250 0.4400 1.2950 0.6500 ;
        RECT 1.9600 0.4300 2.0500 0.6500 ;
        RECT 1.8550 1.2550 2.0550 1.3450 ;
        RECT 1.9550 1.3450 2.0550 1.7200 ;
    END
    ANTENNADIFFAREA 0.375 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2400 0.7950 2.3500 1.1950 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.3500 0.8450 1.6750 0.9450 ;
      RECT 1.5750 0.9450 1.6750 1.1650 ;
      RECT 0.3500 1.3800 0.4500 1.9550 ;
      RECT 0.3500 0.4400 0.4500 0.8450 ;
      RECT 0.3500 1.2800 0.8450 1.3800 ;
      RECT 0.7450 0.9450 0.8450 1.2800 ;
      RECT 1.6800 1.8200 2.3150 1.9200 ;
      RECT 2.2150 1.4900 2.3150 1.8200 ;
      RECT 0.6400 1.4900 1.7800 1.5800 ;
      RECT 1.6800 1.5800 1.7800 1.8200 ;
      RECT 0.6400 1.5800 0.7400 1.9200 ;
      RECT 1.1600 1.5800 1.2600 1.9200 ;
  END
END AOI2XB1_X2M_A12TH

MACRO AOI2XB1_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7800 ;
        RECT 0.6350 0.3200 0.7450 0.6500 ;
        RECT 1.6450 0.3200 1.8150 0.5600 ;
        RECT 2.4700 0.3200 2.6400 0.5600 ;
        RECT 3.0250 0.3200 3.1250 0.6250 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9850 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END A1N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3200 1.2500 2.1950 1.3500 ;
        RECT 1.3200 1.1500 1.4200 1.2500 ;
        RECT 2.0950 0.9450 2.1950 1.2500 ;
        RECT 0.9850 1.0500 1.4200 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.9000 1.7700 1.0000 2.0800 ;
        RECT 1.4200 1.7700 1.5200 2.0800 ;
        RECT 1.9400 1.7700 2.0400 2.0800 ;
        RECT 0.0900 1.6100 0.1900 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1250 0.6500 2.8650 0.7500 ;
        RECT 2.5050 0.7500 2.6050 1.2900 ;
        RECT 2.1650 0.4450 2.3350 0.6500 ;
        RECT 1.1250 0.4400 1.2950 0.6500 ;
        RECT 2.7650 0.4200 2.8650 0.6500 ;
        RECT 2.5050 1.2900 3.1250 1.3900 ;
        RECT 2.5050 1.3900 2.6050 1.7200 ;
        RECT 3.0250 1.3900 3.1250 1.7250 ;
    END
    ANTENNADIFFAREA 0.646875 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7250 0.8500 3.1500 0.9500 ;
    END
    ANTENNAGATEAREA 0.2313 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 1.5400 1.0500 1.9400 1.1500 ;
      RECT 0.3500 0.8500 1.6400 0.9500 ;
      RECT 1.5400 0.9500 1.6400 1.0500 ;
      RECT 0.3500 1.3500 0.4500 1.7800 ;
      RECT 0.3500 0.4650 0.4500 0.8500 ;
      RECT 0.3500 1.2500 0.8400 1.3500 ;
      RECT 0.7400 0.9500 0.8400 1.2500 ;
      RECT 2.2000 1.8200 2.8650 1.9200 ;
      RECT 2.7650 1.4900 2.8650 1.8200 ;
      RECT 0.6400 1.4700 2.3000 1.5700 ;
      RECT 2.2000 1.5700 2.3000 1.8200 ;
      RECT 0.6400 1.5700 0.7400 1.9000 ;
      RECT 1.1600 1.5700 1.2600 1.9000 ;
      RECT 1.6800 1.5700 1.7800 1.9000 ;
  END
END AOI2XB1_X3M_A12TH

MACRO AOI2XB1_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.6500 ;
        RECT 0.6500 0.3200 0.7600 0.6500 ;
        RECT 1.6600 0.3200 1.8300 0.5600 ;
        RECT 2.7050 0.3200 2.8750 0.5600 ;
        RECT 3.2350 0.3200 3.4050 0.5600 ;
        RECT 3.7900 0.3200 3.8900 0.6300 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 1.0500 0.6400 1.1500 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END A1N

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8700 0.8500 3.3100 0.9500 ;
    END
    ANTENNAGATEAREA 0.3084 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.0500 1.4300 1.1550 ;
        RECT 1.3300 1.1550 1.4300 1.2500 ;
        RECT 1.3300 1.2500 2.1500 1.3500 ;
        RECT 2.0500 1.1550 2.1500 1.2500 ;
        RECT 2.0500 1.0550 2.4750 1.1550 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0000 1.2500 3.6350 1.3500 ;
        RECT 3.0000 1.3500 3.1100 1.7200 ;
        RECT 3.5250 1.3500 3.6350 1.7150 ;
        RECT 3.4500 0.7500 3.5500 1.2500 ;
        RECT 1.1400 0.6500 3.6300 0.7500 ;
        RECT 1.1400 0.4400 1.3100 0.6500 ;
        RECT 2.1800 0.4400 2.3500 0.6500 ;
        RECT 3.5300 0.4200 3.6300 0.6500 ;
        RECT 3.0100 0.4150 3.1100 0.6500 ;
    END
    ANTENNADIFFAREA 0.75 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.0950 1.7700 0.1950 2.0800 ;
        RECT 0.9150 1.7700 1.0150 2.0800 ;
        RECT 1.4350 1.7700 1.5350 2.0800 ;
        RECT 1.9550 1.7700 2.0550 2.0800 ;
        RECT 2.4750 1.7700 2.5750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 0.8500 2.7300 0.9500 ;
      RECT 2.6300 0.9500 2.7300 1.1950 ;
      RECT 0.3550 1.4100 0.4550 1.7450 ;
      RECT 0.3550 0.5050 0.4550 0.8500 ;
      RECT 0.3550 1.3100 0.8600 1.4100 ;
      RECT 0.7600 1.1550 0.8600 1.3100 ;
      RECT 0.7600 0.9500 0.8650 1.1550 ;
      RECT 1.5550 0.9500 1.9350 1.0400 ;
      RECT 2.7000 1.8200 3.8900 1.9200 ;
      RECT 3.7900 1.5100 3.8900 1.8200 ;
      RECT 0.6550 1.5100 2.8350 1.6000 ;
      RECT 2.7000 1.6000 2.8350 1.8200 ;
      RECT 3.2650 1.4900 3.3750 1.8200 ;
      RECT 0.6550 1.6000 0.7550 1.9400 ;
      RECT 1.1750 1.6000 1.2750 1.9400 ;
      RECT 1.6950 1.6000 1.7950 1.9400 ;
      RECT 2.2150 1.6000 2.3150 1.9400 ;
  END
END AOI2XB1_X4M_A12TH

MACRO AOI2XB1_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7450 ;
        RECT 0.6150 0.3200 0.7150 0.7400 ;
        RECT 0.9100 0.3200 1.0200 0.6500 ;
        RECT 1.9200 0.3200 2.0900 0.5400 ;
        RECT 2.9600 0.3200 3.1300 0.5400 ;
        RECT 4.0050 0.3200 4.1750 0.5550 ;
        RECT 4.5350 0.3200 4.7050 0.7400 ;
        RECT 5.0550 0.3200 5.2250 0.7400 ;
        RECT 5.6100 0.3200 5.7100 0.8350 ;
    END
  END VSS

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1650 1.0500 0.6050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1482 ;
  END A1N

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2100 1.0500 4.9200 1.1500 ;
    END
    ANTENNAGATEAREA 0.4626 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 1.2500 3.4500 1.3500 ;
        RECT 3.3500 1.1550 3.4500 1.2500 ;
        RECT 1.6000 1.1500 1.7000 1.2500 ;
        RECT 2.3350 1.0600 2.7150 1.2500 ;
        RECT 3.3500 1.0550 3.7750 1.1550 ;
        RECT 1.2500 1.0500 1.7000 1.1500 ;
    END
    ANTENNAGATEAREA 0.54 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3000 1.2500 5.4500 1.3500 ;
        RECT 4.3000 1.3500 4.4100 1.7200 ;
        RECT 4.8300 1.3500 4.9300 1.7200 ;
        RECT 5.3500 1.3500 5.4500 1.7200 ;
        RECT 5.0500 0.9500 5.1500 1.2500 ;
        RECT 4.3100 0.8500 5.4500 0.9500 ;
        RECT 4.3100 0.7550 4.4100 0.8500 ;
        RECT 4.8300 0.4400 4.9300 0.8500 ;
        RECT 5.3500 0.4400 5.4500 0.8500 ;
        RECT 1.4000 0.6550 4.4100 0.7550 ;
        RECT 3.4800 0.4650 3.6500 0.6550 ;
        RECT 4.3100 0.4400 4.4100 0.6550 ;
        RECT 1.4000 0.4200 1.5700 0.6550 ;
        RECT 2.4400 0.4200 2.6100 0.6550 ;
    END
    ANTENNADIFFAREA 1.125 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 1.1750 1.7700 1.2750 2.0800 ;
        RECT 1.6950 1.7700 1.7950 2.0800 ;
        RECT 2.2150 1.7700 2.3150 2.0800 ;
        RECT 2.7350 1.7700 2.8350 2.0800 ;
        RECT 3.2550 1.7700 3.3550 2.0800 ;
        RECT 3.7750 1.7700 3.8750 2.0800 ;
        RECT 0.0950 1.7100 0.1950 2.0800 ;
        RECT 0.6150 1.7000 0.7150 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 0.4250 0.4550 0.8600 ;
      RECT 0.3550 0.8600 4.0300 0.9600 ;
      RECT 0.3600 1.2900 1.1200 1.3900 ;
      RECT 0.3600 1.3900 0.4600 1.8700 ;
      RECT 1.0200 0.9600 1.1200 1.2900 ;
      RECT 3.9300 0.9600 4.0300 1.1800 ;
      RECT 1.8150 0.8600 2.1950 1.1000 ;
      RECT 2.8550 0.8600 3.2350 1.1000 ;
      RECT 4.0250 1.8200 5.7100 1.9200 ;
      RECT 5.6100 1.5100 5.7100 1.8200 ;
      RECT 0.9150 1.5100 4.1600 1.6000 ;
      RECT 4.0250 1.6000 4.1600 1.8200 ;
      RECT 4.5650 1.4900 4.6750 1.8200 ;
      RECT 5.0850 1.4900 5.1950 1.8200 ;
      RECT 0.9150 1.6000 1.0150 1.9400 ;
      RECT 1.4350 1.6000 1.5350 1.9400 ;
      RECT 1.9550 1.6000 2.0550 1.9400 ;
      RECT 2.4750 1.6000 2.5750 1.9400 ;
      RECT 2.9950 1.6000 3.0950 1.9400 ;
      RECT 3.5150 1.6000 3.6150 1.9400 ;
  END
END AOI2XB1_X6M_A12TH

MACRO AOI2XB1_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7500 ;
        RECT 0.6100 0.3200 0.7100 0.7500 ;
        RECT 0.8800 0.3200 0.9900 0.6500 ;
        RECT 1.8700 0.3200 2.0800 0.4100 ;
        RECT 2.9100 0.3200 3.1200 0.4100 ;
        RECT 3.9500 0.3200 4.1600 0.4100 ;
        RECT 5.0300 0.3200 5.2400 0.4100 ;
        RECT 5.6550 0.3200 5.7550 0.4300 ;
        RECT 6.1750 0.3200 6.2750 0.4300 ;
        RECT 6.6950 0.3200 6.7950 0.4300 ;
        RECT 7.2150 0.3200 7.3150 0.6250 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2700 0.8500 6.1900 0.9500 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5650 1.2500 4.4700 1.3500 ;
        RECT 1.5650 1.1550 1.6650 1.2500 ;
        RECT 4.3700 1.1500 4.4700 1.2500 ;
        RECT 2.3100 1.0600 2.6800 1.2500 ;
        RECT 3.3500 1.0600 3.7200 1.2500 ;
        RECT 1.2550 1.0550 1.6650 1.1550 ;
        RECT 4.3700 1.0600 4.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.72 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3700 0.5700 7.0900 0.7500 ;
        RECT 6.6100 0.7500 6.7900 1.2100 ;
        RECT 5.3600 0.4600 5.5300 0.5700 ;
        RECT 5.8800 0.4600 6.0500 0.5700 ;
        RECT 6.4000 0.4600 6.5700 0.5700 ;
        RECT 6.9200 0.4600 7.0900 0.5700 ;
        RECT 1.3700 0.4400 1.5400 0.5700 ;
        RECT 2.4100 0.4400 2.5800 0.5700 ;
        RECT 3.4500 0.4400 3.6200 0.5700 ;
        RECT 4.4900 0.4400 4.6600 0.5700 ;
        RECT 5.3850 1.2100 7.0600 1.3900 ;
        RECT 5.3850 1.3900 5.4950 1.7200 ;
        RECT 5.9100 1.3900 6.0200 1.7200 ;
        RECT 6.4300 1.3900 6.5400 1.7200 ;
        RECT 6.9500 1.3900 7.0600 1.7200 ;
    END
    ANTENNADIFFAREA 1.5 ;
  END Y

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.0500 0.7600 1.1500 ;
    END
    ANTENNAGATEAREA 0.195 ;
  END A1N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1450 1.7700 1.2450 2.0800 ;
        RECT 1.6650 1.7700 1.7650 2.0800 ;
        RECT 2.1850 1.7700 2.2850 2.0800 ;
        RECT 2.7050 1.7700 2.8050 2.0800 ;
        RECT 3.2250 1.7700 3.3250 2.0800 ;
        RECT 3.7450 1.7700 3.8450 2.0800 ;
        RECT 4.2650 1.7700 4.3650 2.0800 ;
        RECT 4.7900 1.7700 4.8900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 5.0750 1.8200 7.3200 1.9200 ;
      RECT 7.2100 1.4900 7.3200 1.8200 ;
      RECT 0.8850 1.5100 5.2100 1.6000 ;
      RECT 5.0750 1.6000 5.2100 1.8200 ;
      RECT 5.6500 1.4900 5.7600 1.8200 ;
      RECT 6.1700 1.4900 6.2800 1.8200 ;
      RECT 6.6900 1.4900 6.8000 1.8200 ;
      RECT 0.8850 1.6000 0.9850 1.9400 ;
      RECT 1.4050 1.6000 1.5050 1.9400 ;
      RECT 1.9250 1.6000 2.0250 1.9400 ;
      RECT 2.4450 1.6000 2.5450 1.9400 ;
      RECT 2.9650 1.6000 3.0650 1.9400 ;
      RECT 3.4850 1.6000 3.5850 1.9400 ;
      RECT 4.0050 1.6000 4.1050 1.9400 ;
      RECT 4.5250 1.6000 4.6250 1.9400 ;
      RECT 0.3500 0.4850 0.4500 0.8600 ;
      RECT 0.3500 1.3900 0.4500 1.7200 ;
      RECT 0.3500 0.8600 5.0750 0.9600 ;
      RECT 0.3500 1.2900 1.0900 1.3900 ;
      RECT 0.9900 0.9600 1.0950 1.1200 ;
      RECT 0.9900 1.1200 1.0900 1.2900 ;
      RECT 4.9750 0.9600 5.0750 1.2250 ;
      RECT 1.7950 0.8600 2.1650 1.0950 ;
      RECT 2.8300 0.8600 3.2000 1.0950 ;
      RECT 3.8700 0.8600 4.2400 1.0950 ;
  END
END AOI2XB1_X8M_A12TH

MACRO AOI31_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1250 0.3200 0.2250 0.7150 ;
        RECT 1.2000 0.3200 1.3000 0.5050 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.5650 ;
        RECT 1.2000 1.5650 1.3500 1.6550 ;
        RECT 0.8300 0.6000 1.3500 0.7000 ;
        RECT 1.2000 1.6550 1.3000 1.9900 ;
        RECT 0.8300 0.4100 1.0000 0.6000 ;
    END
    ANTENNADIFFAREA 0.160125 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 0.8500 0.9100 0.9500 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.2500 0.7100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 0.8100 0.3500 0.9200 ;
        RECT 0.2500 0.9200 0.3500 1.1300 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6650 1.6250 0.7650 2.0800 ;
        RECT 0.1250 1.5750 0.2250 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8900 1.1500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0363 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.3900 1.4450 1.0300 1.5350 ;
      RECT 0.9400 1.5350 1.0300 1.9900 ;
      RECT 0.3900 1.5350 0.4800 1.9900 ;
  END
END AOI31_X0P5M_A12TH

MACRO AOI31_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.1000 0.3200 0.2000 0.6300 ;
        RECT 1.2000 0.3200 1.3000 0.4400 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2900 1.2500 0.7100 1.3500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7450 1.3500 1.5350 ;
        RECT 1.2000 1.5350 1.3500 1.6250 ;
        RECT 0.7950 0.6450 1.3500 0.7450 ;
        RECT 1.2000 1.6250 1.3000 1.9650 ;
        RECT 0.7950 0.4200 0.9650 0.6450 ;
    END
    ANTENNADIFFAREA 0.235875 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 0.8500 0.9100 0.9500 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A0

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1450 0.7800 0.3500 1.1050 ;
    END
    ANTENNAGATEAREA 0.0693 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1000 1.7150 0.2000 2.0800 ;
        RECT 0.6500 1.7150 0.7500 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.8850 1.1500 1.3050 ;
    END
    ANTENNAGATEAREA 0.0516 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.3650 1.5150 1.0350 1.6050 ;
      RECT 0.9450 1.6050 1.0350 1.9650 ;
      RECT 0.3650 1.6050 0.4550 1.9650 ;
  END
END AOI31_X0P7M_A12TH

MACRO AOI31_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 1.2100 0.3200 1.3100 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7400 1.3500 1.5000 ;
        RECT 1.2100 1.5000 1.3500 1.6000 ;
        RECT 0.8300 0.6400 1.3500 0.7400 ;
        RECT 1.2100 1.6000 1.3100 1.9150 ;
        RECT 0.8300 0.4350 1.0000 0.6400 ;
    END
    ANTENNADIFFAREA 0.3243 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2500 0.9500 1.4000 ;
        RECT 0.7600 1.0800 0.9500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2850 1.2500 0.5900 1.3500 ;
        RECT 0.4900 1.0800 0.5900 1.2500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0200 0.3900 1.1500 ;
    END
    ANTENNAGATEAREA 0.0978 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6450 1.7700 0.7450 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8850 1.1500 1.3150 ;
    END
    ANTENNAGATEAREA 0.0729 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.3800 1.5150 1.0500 1.6050 ;
      RECT 0.9500 1.6050 1.0500 1.9450 ;
      RECT 0.3800 1.6050 0.4800 1.9450 ;
  END
END AOI31_X1M_A12TH

MACRO AOI31_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.3150 0.3200 0.4850 0.5650 ;
        RECT 2.1900 0.3200 2.2900 0.6850 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.7850 1.7500 1.3150 ;
        RECT 1.6500 1.3150 2.0300 1.4150 ;
        RECT 1.3750 0.6850 2.0300 0.7850 ;
        RECT 1.9300 1.4150 2.0300 1.7200 ;
        RECT 1.3750 0.6700 1.5700 0.6850 ;
        RECT 1.9300 0.4150 2.0300 0.6850 ;
    END
    ANTENNADIFFAREA 0.32255 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2550 1.0050 1.5500 1.1050 ;
        RECT 1.4500 1.1050 1.5500 1.3050 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6800 1.2500 1.1100 1.3500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 1.0500 0.5100 1.1500 ;
    END
    ANTENNAGATEAREA 0.1386 ;
  END A2

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8850 1.0500 2.3150 1.1500 ;
    END
    ANTENNAGATEAREA 0.1032 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3500 1.7150 0.4500 2.0800 ;
        RECT 0.8700 1.7150 0.9700 2.0800 ;
        RECT 1.3900 1.7150 1.4900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 0.6850 1.2650 0.7850 ;
      RECT 1.0750 0.6700 1.2650 0.6850 ;
      RECT 0.6150 0.4150 0.7050 0.6850 ;
      RECT 0.0950 0.4150 0.1850 0.6850 ;
      RECT 0.8150 0.4850 1.8200 0.5750 ;
      RECT 1.6700 1.8200 2.2900 1.9200 ;
      RECT 2.1900 1.5100 2.2900 1.8200 ;
      RECT 0.0900 1.5200 1.7700 1.6100 ;
      RECT 1.6700 1.6100 1.7700 1.8200 ;
      RECT 0.0900 1.6100 0.1900 1.9450 ;
      RECT 0.6100 1.6100 0.7100 1.9450 ;
      RECT 1.1300 1.6100 1.2300 1.9450 ;
  END
END AOI31_X1P4M_A12TH

MACRO AOI31_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.6300 0.3200 0.7300 0.6950 ;
        RECT 2.2000 0.3200 2.3000 0.6350 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.2500 1.9350 1.3500 ;
        RECT 1.0400 1.0400 1.1400 1.2500 ;
        RECT 1.8350 1.0400 1.9350 1.2500 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8050 1.4500 2.1250 1.5500 ;
        RECT 2.0250 1.1950 2.1250 1.4500 ;
        RECT 0.8050 1.0600 0.9050 1.4500 ;
        RECT 2.0250 1.0950 2.2550 1.1950 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A2

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0500 1.6600 1.1600 ;
    END
    ANTENNAGATEAREA 0.1956 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.4900 1.1600 ;
    END
    ANTENNAGATEAREA 0.1458 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3550 0.8500 0.9500 0.9500 ;
        RECT 0.6000 0.9500 0.7000 1.2500 ;
        RECT 0.8500 0.5800 0.9500 0.8500 ;
        RECT 0.3550 0.5250 0.4550 0.8500 ;
        RECT 0.3550 1.2500 0.7000 1.3500 ;
        RECT 0.8500 0.4800 1.5200 0.5800 ;
        RECT 0.3550 1.3500 0.4550 1.7350 ;
        RECT 1.4200 0.5800 1.5200 0.9000 ;
    END
    ANTENNADIFFAREA 0.47155 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.8900 1.8200 0.9900 2.0800 ;
        RECT 1.4200 1.8200 1.5200 2.0800 ;
        RECT 1.9400 1.8200 2.0400 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.6250 1.6400 2.3050 1.7300 ;
      RECT 2.2150 1.3400 2.3050 1.6400 ;
      RECT 0.1000 1.8300 0.7150 1.9200 ;
      RECT 0.6250 1.7300 0.7150 1.8300 ;
      RECT 0.6250 1.5000 0.7150 1.6400 ;
      RECT 0.1000 1.4900 0.1900 1.8300 ;
      RECT 1.1250 1.7300 1.2950 1.9300 ;
      RECT 1.6450 1.7300 1.8150 1.9300 ;
  END
END AOI31_X2M_A12TH

MACRO AOI31_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0850 0.3200 0.1950 0.6300 ;
        RECT 0.6050 0.3200 0.7150 0.6300 ;
        RECT 2.6550 0.3200 2.8250 0.5400 ;
        RECT 3.2100 0.3200 3.3100 0.7750 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.7800 2.5500 1.3000 ;
        RECT 2.4500 1.3000 3.3100 1.4000 ;
        RECT 1.9100 0.7600 2.5500 0.7800 ;
        RECT 2.6900 1.4000 2.7900 1.7200 ;
        RECT 3.2100 1.4000 3.3100 1.7700 ;
        RECT 1.9100 0.7800 2.0100 0.8700 ;
        RECT 1.9100 0.6600 3.0850 0.7600 ;
        RECT 2.9150 0.4350 3.0850 0.6600 ;
        RECT 2.4300 0.4100 2.5300 0.6600 ;
    END
    ANTENNADIFFAREA 0.666225 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8550 1.0500 2.3250 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0550 1.0500 1.5200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.0350 0.7500 1.1500 ;
    END
    ANTENNAGATEAREA 0.2934 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 0.6100 1.7700 0.7100 2.0800 ;
        RECT 1.1300 1.7700 1.2300 2.0800 ;
        RECT 1.6500 1.7700 1.7500 2.0800 ;
        RECT 2.1700 1.7700 2.2700 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6950 1.0200 3.1050 1.1550 ;
    END
    ANTENNAGATEAREA 0.2187 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 2.4300 1.8200 3.0500 1.9200 ;
      RECT 2.9500 1.5100 3.0500 1.8200 ;
      RECT 0.3500 1.5000 2.5300 1.5900 ;
      RECT 2.4300 1.5900 2.5300 1.8200 ;
      RECT 0.3500 1.5900 0.4500 1.9200 ;
      RECT 0.8700 1.5900 0.9700 1.9200 ;
      RECT 1.3900 1.5900 1.4900 1.9200 ;
      RECT 1.9100 1.5900 2.0100 1.9200 ;
      RECT 0.3550 0.8100 1.4850 0.9000 ;
      RECT 1.3950 0.7100 1.4850 0.8100 ;
      RECT 0.8750 0.4400 0.9650 0.8100 ;
      RECT 0.3550 0.4400 0.4450 0.8100 ;
      RECT 1.1350 0.4800 2.3050 0.5700 ;
      RECT 1.1350 0.5700 1.2250 0.6900 ;
      RECT 1.6500 0.5700 1.7500 0.8900 ;
  END
END AOI31_X3M_A12TH

MACRO AOI21B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7300 ;
        RECT 1.1300 0.3200 1.2300 0.7000 ;
        RECT 1.7100 0.3200 1.8100 0.6900 ;
        RECT 2.2200 0.3200 2.3200 0.7600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.4600 1.5500 0.8000 ;
        RECT 0.6100 0.8000 1.5500 0.9000 ;
        RECT 1.2500 0.9000 1.3500 1.2650 ;
        RECT 0.6100 0.4550 0.7100 0.8000 ;
        RECT 1.2500 1.2650 1.4900 1.3650 ;
        RECT 1.3900 1.3650 1.4900 1.7200 ;
    END
    ANTENNADIFFAREA 0.375 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 2.2250 1.5000 2.3250 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9000 0.1600 1.2500 ;
        RECT 0.0500 1.2500 1.1500 1.3500 ;
        RECT 1.0250 1.0100 1.1500 1.2500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0500 0.8650 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9000 1.0500 2.3300 1.1500 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END B0N
  OBS
    LAYER M1 ;
      RECT 1.1300 1.8200 1.7500 1.9200 ;
      RECT 1.6500 1.4900 1.7500 1.8200 ;
      RECT 0.0900 1.4800 1.2300 1.5900 ;
      RECT 1.1300 1.5900 1.2300 1.8200 ;
      RECT 0.0900 1.5900 0.1900 1.9100 ;
      RECT 0.6100 1.5900 0.7100 1.9100 ;
      RECT 1.9600 1.3800 2.0600 1.9500 ;
      RECT 1.6650 1.2800 2.0600 1.3800 ;
      RECT 1.6650 0.8100 2.0600 0.9100 ;
      RECT 1.9600 0.6550 2.0600 0.8100 ;
      RECT 1.6650 1.1800 1.7650 1.2800 ;
      RECT 1.5300 1.0800 1.7650 1.1800 ;
      RECT 1.6650 0.9100 1.7650 1.0800 ;
  END
END AOI21B_X2M_A12TH

MACRO AOI21B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7300 ;
        RECT 1.1300 0.3200 1.2300 0.5100 ;
        RECT 1.9550 0.3200 2.0550 0.5100 ;
        RECT 2.4750 0.3200 2.5750 0.7100 ;
        RECT 3.0100 0.3200 3.1100 0.8400 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5750 0.6500 2.3150 0.7500 ;
        RECT 1.9250 0.7500 2.0250 1.2500 ;
        RECT 1.6500 0.4750 1.7500 0.6500 ;
        RECT 2.2150 0.4750 2.3150 0.6500 ;
        RECT 0.5750 0.4200 0.7450 0.6500 ;
        RECT 1.9250 1.2500 2.5450 1.3500 ;
        RECT 1.9250 1.3500 2.0250 1.7200 ;
        RECT 2.4450 1.3500 2.5450 1.7200 ;
    END
    ANTENNADIFFAREA 0.6396 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 1.3900 1.7700 1.4900 2.0800 ;
        RECT 3.0150 1.6850 3.1150 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9000 0.3500 1.2500 ;
        RECT 0.2500 1.2500 1.0900 1.3500 ;
        RECT 0.9900 1.1700 1.0900 1.2500 ;
        RECT 0.9900 1.0600 1.3600 1.1700 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9500 1.5900 1.2900 ;
        RECT 0.7700 0.8500 1.5900 0.9500 ;
        RECT 0.7700 0.9500 0.8700 1.0500 ;
        RECT 0.4700 1.0500 0.8700 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0400 1.0100 3.1500 1.4250 ;
    END
    ANTENNAGATEAREA 0.0648 ;
  END B0N
  OBS
    LAYER M1 ;
      RECT 1.6600 1.8300 2.2850 1.9200 ;
      RECT 2.1850 1.5100 2.2850 1.8300 ;
      RECT 0.0900 1.4800 1.7600 1.5900 ;
      RECT 1.6600 1.5900 1.7600 1.8300 ;
      RECT 0.0900 1.5900 0.1900 1.9100 ;
      RECT 0.6100 1.5900 0.7100 1.9100 ;
      RECT 1.1300 1.5900 1.2300 1.9100 ;
      RECT 2.7500 1.5550 2.8500 1.9400 ;
      RECT 2.6500 1.4550 2.8500 1.5550 ;
      RECT 2.6500 1.1600 2.7500 1.4550 ;
      RECT 2.1500 1.0500 2.7500 1.1600 ;
      RECT 2.6500 0.9350 2.7500 1.0500 ;
      RECT 2.6500 0.8350 2.8500 0.9350 ;
      RECT 2.7500 0.4850 2.8500 0.8350 ;
  END
END AOI21B_X3M_A12TH

MACRO AOI21B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7300 ;
        RECT 1.0750 0.3200 1.2850 0.4500 ;
        RECT 2.1700 0.3200 2.2700 0.6750 ;
        RECT 2.7450 0.3200 2.8450 0.5100 ;
        RECT 3.2650 0.3200 3.3650 0.6900 ;
        RECT 3.7900 0.3200 3.8900 0.7450 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7650 0.8500 1.5800 0.9500 ;
        RECT 1.4800 0.9500 1.5800 1.0350 ;
        RECT 0.7650 0.9500 0.8650 1.0250 ;
        RECT 1.4800 1.0350 1.9100 1.1350 ;
        RECT 0.4700 1.0250 0.8650 1.1250 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 2.1500 1.3500 ;
        RECT 0.9900 1.0600 1.3700 1.2500 ;
        RECT 2.0200 1.0200 2.1500 1.2500 ;
        RECT 0.2500 0.9950 0.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4100 1.0500 3.8400 1.1500 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END B0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 1.2500 3.0500 1.3500 ;
        RECT 2.4300 1.3500 2.5300 1.7200 ;
        RECT 2.9500 1.3500 3.0500 1.7200 ;
        RECT 2.2500 0.9000 2.3500 1.2500 ;
        RECT 1.6850 0.8000 3.1050 0.9000 ;
        RECT 1.6850 0.7300 1.7850 0.8000 ;
        RECT 2.4850 0.4650 2.5850 0.8000 ;
        RECT 3.0050 0.4650 3.1050 0.8000 ;
        RECT 0.5750 0.6300 1.7850 0.7300 ;
        RECT 0.5750 0.4400 0.7450 0.6300 ;
        RECT 1.6150 0.4400 1.7850 0.6300 ;
    END
    ANTENNADIFFAREA 0.75 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 1.3900 1.7700 1.4900 2.0800 ;
        RECT 1.9100 1.7650 2.0100 2.0800 ;
        RECT 3.7950 1.6850 3.8950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1700 1.8300 3.3100 1.9200 ;
      RECT 3.2100 1.5100 3.3100 1.8300 ;
      RECT 0.0900 1.5200 2.2700 1.6200 ;
      RECT 2.1700 1.6200 2.2700 1.8300 ;
      RECT 2.6900 1.5000 2.7900 1.8300 ;
      RECT 0.0900 1.6200 0.1900 1.9500 ;
      RECT 0.6100 1.6200 0.7100 1.9600 ;
      RECT 1.1300 1.6200 1.2300 1.9550 ;
      RECT 1.6500 1.6200 1.7500 1.9600 ;
      RECT 3.5300 1.3750 3.6300 1.7400 ;
      RECT 3.2050 1.2750 3.6300 1.3750 ;
      RECT 3.2050 0.8400 3.6300 0.9400 ;
      RECT 3.5300 0.5100 3.6300 0.8400 ;
      RECT 3.2050 1.1300 3.3050 1.2750 ;
      RECT 2.8150 1.0300 3.3050 1.1300 ;
      RECT 3.2050 0.9400 3.3050 1.0300 ;
  END
END AOI21B_X4M_A12TH

MACRO AOI21B_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7200 ;
        RECT 1.1250 0.3200 1.2350 0.5100 ;
        RECT 2.1650 0.3200 2.2750 0.5100 ;
        RECT 3.2100 0.3200 3.3100 0.6850 ;
        RECT 3.7650 0.3200 3.8750 0.6950 ;
        RECT 4.2850 0.3200 4.3950 0.6950 ;
        RECT 4.8100 0.3200 4.9100 0.9050 ;
        RECT 5.0900 0.3200 5.1900 0.7150 ;
        RECT 5.6100 0.3200 5.7100 0.7350 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9800 0.3500 1.2500 ;
        RECT 0.2500 1.2500 3.2050 1.3500 ;
        RECT 0.9900 1.0600 1.3700 1.2500 ;
        RECT 2.0300 1.0600 2.4100 1.2500 ;
        RECT 3.1050 1.0150 3.2050 1.2500 ;
    END
    ANTENNAGATEAREA 0.54 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2500 1.0350 5.6000 1.2150 ;
    END
    ANTENNAGATEAREA 0.129 ;
  END B0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5100 1.2500 4.6500 1.3500 ;
        RECT 3.5100 1.3500 3.6100 1.7100 ;
        RECT 4.0300 1.3500 4.1300 1.7100 ;
        RECT 4.5500 1.3500 4.6500 1.7100 ;
        RECT 3.5100 0.8950 3.6100 1.2500 ;
        RECT 2.7250 0.7950 4.6500 0.8950 ;
        RECT 2.7250 0.7300 2.8250 0.7950 ;
        RECT 3.5100 0.5000 3.6100 0.7950 ;
        RECT 4.0300 0.5000 4.1300 0.7950 ;
        RECT 4.5500 0.5000 4.6500 0.7950 ;
        RECT 0.5750 0.6300 2.8250 0.7300 ;
        RECT 0.5750 0.4350 0.7450 0.6300 ;
        RECT 1.6150 0.4350 1.7850 0.6300 ;
        RECT 2.6550 0.4350 2.8250 0.6300 ;
    END
    ANTENNADIFFAREA 1.125 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 0.8500 2.6200 0.9500 ;
        RECT 0.7700 0.9500 0.8700 1.0500 ;
        RECT 1.5100 0.9500 1.8900 1.1200 ;
        RECT 2.5200 0.9500 2.6200 1.0500 ;
        RECT 0.4700 1.0500 0.8700 1.1500 ;
        RECT 2.5200 1.0500 2.9500 1.1500 ;
    END
    ANTENNAGATEAREA 0.54 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 1.3900 1.7700 1.4900 2.0800 ;
        RECT 2.4300 1.7700 2.5300 2.0800 ;
        RECT 2.9500 1.7700 3.0500 2.0800 ;
        RECT 1.9100 1.7650 2.0100 2.0800 ;
        RECT 5.0900 1.6800 5.1900 2.0800 ;
        RECT 5.6100 1.6700 5.7100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.2350 1.8300 4.9100 1.9200 ;
      RECT 4.8100 1.4900 4.9100 1.8300 ;
      RECT 0.0900 1.4700 3.3350 1.5700 ;
      RECT 3.2350 1.5700 3.3350 1.8300 ;
      RECT 3.7700 1.4850 3.8700 1.8300 ;
      RECT 4.2900 1.4900 4.3900 1.8300 ;
      RECT 0.0900 1.5700 0.1900 1.9000 ;
      RECT 0.6100 1.5700 0.7100 1.9000 ;
      RECT 1.1300 1.5700 1.2300 1.9000 ;
      RECT 1.6500 1.5700 1.7500 1.9050 ;
      RECT 2.1700 1.5700 2.2700 1.9000 ;
      RECT 2.6900 1.5700 2.7900 1.9050 ;
      RECT 5.3500 1.5800 5.4500 1.9300 ;
      RECT 5.0200 1.4800 5.4500 1.5800 ;
      RECT 5.0200 0.8250 5.4500 0.9250 ;
      RECT 5.3500 0.4100 5.4500 0.8250 ;
      RECT 5.0200 1.1250 5.1200 1.4800 ;
      RECT 3.7900 1.0250 5.1200 1.1250 ;
      RECT 5.0200 0.9250 5.1200 1.0250 ;
  END
END AOI21B_X6M_A12TH

MACRO AOI21B_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6450 ;
        RECT 1.1300 0.3200 1.2300 0.4300 ;
        RECT 2.1700 0.3200 2.2700 0.4300 ;
        RECT 3.2100 0.3200 3.3100 0.4300 ;
        RECT 4.2700 0.3200 4.3700 0.4300 ;
        RECT 4.7900 0.3200 4.8900 0.4300 ;
        RECT 5.3100 0.3200 5.4100 0.4300 ;
        RECT 5.8300 0.3200 5.9300 0.4300 ;
        RECT 6.3500 0.3200 6.4500 0.6050 ;
        RECT 6.6400 0.3200 6.7400 0.6100 ;
        RECT 7.1600 0.3200 7.2600 0.6100 ;
    END
  END VSS

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.7650 1.0400 7.1500 1.1500 ;
    END
    ANTENNAGATEAREA 0.1704 ;
  END B0N

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9200 0.3500 1.2500 ;
        RECT 0.2500 1.2500 4.1900 1.3500 ;
        RECT 0.9900 1.0600 1.3700 1.2500 ;
        RECT 2.0250 1.0600 2.4100 1.2500 ;
        RECT 3.0650 1.0600 3.4500 1.2500 ;
        RECT 4.0900 0.9450 4.1900 1.2500 ;
    END
    ANTENNAGATEAREA 0.72 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.4450 2.7200 ;
        RECT 2.9500 1.7700 3.0500 2.0800 ;
        RECT 3.4700 1.7700 3.5700 2.0800 ;
        RECT 3.9900 1.7700 4.0900 2.0800 ;
        RECT 0.3500 1.7600 0.4500 2.0800 ;
        RECT 0.8700 1.7600 0.9700 2.0800 ;
        RECT 1.3900 1.7600 1.4900 2.0800 ;
        RECT 2.4300 1.7600 2.5300 2.0800 ;
        RECT 1.9100 1.7550 2.0100 2.0800 ;
        RECT 6.6400 1.6900 6.7400 2.0800 ;
        RECT 7.1600 1.6900 7.2600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6100 0.7900 4.7900 1.2000 ;
        RECT 4.5300 1.2000 6.1900 1.3800 ;
        RECT 3.7950 0.7300 6.2050 0.7900 ;
        RECT 4.5300 1.3800 4.6300 1.7250 ;
        RECT 5.0500 1.3800 5.1500 1.7200 ;
        RECT 5.5700 1.3800 5.6700 1.7200 ;
        RECT 6.0900 1.3800 6.1900 1.7200 ;
        RECT 0.5750 0.6100 6.2050 0.7300 ;
        RECT 0.5750 0.5500 3.9750 0.6100 ;
        RECT 4.5200 0.4150 4.6400 0.6100 ;
        RECT 5.0400 0.4150 5.1600 0.6100 ;
        RECT 5.5600 0.4150 5.6800 0.6100 ;
        RECT 6.0850 0.4150 6.2050 0.6100 ;
        RECT 0.5750 0.4200 0.7450 0.5500 ;
        RECT 1.6150 0.4200 1.7850 0.5500 ;
        RECT 2.6550 0.4200 2.8250 0.5500 ;
        RECT 3.6950 0.4200 3.8650 0.5500 ;
    END
    ANTENNADIFFAREA 1.5 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 0.8500 3.6850 0.9500 ;
        RECT 0.7700 0.9500 0.8700 1.0500 ;
        RECT 1.5100 0.9500 1.8900 1.0950 ;
        RECT 2.5500 0.9500 2.9300 1.0950 ;
        RECT 3.5850 0.9500 3.6850 1.0250 ;
        RECT 0.4700 1.0500 0.8700 1.1500 ;
        RECT 3.5850 1.0250 3.9800 1.1250 ;
    END
    ANTENNAGATEAREA 0.72 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 4.2600 1.8300 6.4500 1.9200 ;
      RECT 6.3500 1.4900 6.4500 1.8300 ;
      RECT 0.0900 1.4700 4.3600 1.5700 ;
      RECT 4.2600 1.5700 4.3600 1.8300 ;
      RECT 0.0900 1.5700 0.1900 1.9000 ;
      RECT 0.6100 1.5700 0.7100 1.9000 ;
      RECT 1.1300 1.5700 1.2300 1.9000 ;
      RECT 1.6500 1.5700 1.7500 1.9050 ;
      RECT 2.1700 1.5700 2.2700 1.9000 ;
      RECT 2.6900 1.5700 2.7900 1.9050 ;
      RECT 3.2100 1.5700 3.3100 1.9000 ;
      RECT 3.7300 1.5700 3.8300 1.9050 ;
      RECT 4.7900 1.5000 4.8900 1.8300 ;
      RECT 5.3100 1.5100 5.4100 1.8300 ;
      RECT 5.8300 1.5100 5.9300 1.8300 ;
      RECT 6.9000 1.3800 7.0000 1.7450 ;
      RECT 6.4500 1.2800 7.0000 1.3800 ;
      RECT 6.4500 0.7250 7.0000 0.8250 ;
      RECT 6.9000 0.4150 7.0000 0.7250 ;
      RECT 6.4500 1.0200 6.5500 1.2800 ;
      RECT 4.9550 0.9200 6.5500 1.0200 ;
      RECT 6.4500 0.8250 6.5500 0.9200 ;
  END
END AOI21B_X8M_A12TH

MACRO AOI21_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.1150 0.3200 0.2250 0.6700 ;
        RECT 0.9850 0.3200 1.0950 0.6600 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8600 1.1500 1.5050 ;
        RECT 0.9800 1.5050 1.1500 1.8950 ;
        RECT 0.6800 0.7600 1.1500 0.8600 ;
        RECT 0.6800 0.4600 0.7800 0.7600 ;
    END
    ANTENNADIFFAREA 0.189475 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.9600 0.9500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0384 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7300 0.5600 1.1550 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7700 0.1600 1.1600 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3750 1.7250 0.4850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5000 0.7600 1.6000 ;
      RECT 0.6600 1.6000 0.7600 1.9100 ;
      RECT 0.1200 1.6000 0.2200 1.9100 ;
  END
END AOI21_X0P5M_A12TH

MACRO AOI21_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0850 0.3200 0.2550 0.7200 ;
        RECT 0.9850 0.3200 1.0950 0.6000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8050 1.1500 1.5000 ;
        RECT 0.9800 1.5000 1.1500 1.9100 ;
        RECT 0.6500 0.7050 1.1500 0.8050 ;
        RECT 0.6500 0.4300 0.7500 0.7050 ;
    END
    ANTENNADIFFAREA 0.262 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.9250 0.9500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0546 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7300 0.5600 1.1200 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8950 0.1600 1.3050 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3750 1.6900 0.4850 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5000 0.7600 1.6000 ;
      RECT 0.6600 1.6000 0.7600 1.9100 ;
      RECT 0.1200 1.6000 0.2200 1.9100 ;
  END
END AOI21_X0P7M_A12TH

MACRO AOI21_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.0850 0.3200 0.2550 0.5200 ;
        RECT 0.9900 0.3200 1.0900 0.4300 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.6950 0.1600 1.1150 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7200 1.1500 1.5000 ;
        RECT 0.9800 1.5000 1.1500 1.9100 ;
        RECT 0.6050 0.6200 1.1500 0.7200 ;
        RECT 0.6050 0.4100 0.7750 0.6200 ;
    END
    ANTENNADIFFAREA 0.3249 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 0.8900 0.9500 1.3100 ;
    END
    ANTENNAGATEAREA 0.0771 ;
  END B0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.3800 1.7700 0.4800 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8100 0.7250 0.9150 ;
        RECT 0.4500 0.9150 0.5600 1.1200 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5000 0.7600 1.6000 ;
      RECT 0.6600 1.6000 0.7600 1.9100 ;
      RECT 0.1200 1.6000 0.2200 1.9100 ;
  END
END AOI21_X1M_A12TH

MACRO AOI21_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.8700 ;
        RECT 1.2000 0.3200 1.3000 0.6700 ;
        RECT 1.7600 0.3200 1.8600 0.6700 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.3800 1.7400 0.4800 2.0800 ;
        RECT 0.9000 1.7400 1.0000 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.0000 1.7600 1.3850 ;
    END
    ANTENNAGATEAREA 0.1092 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0800 1.2500 1.1600 1.3500 ;
        RECT 1.0700 1.3500 1.1600 1.4200 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9000 1.5500 1.5650 ;
        RECT 1.4500 1.5650 1.6350 1.6550 ;
        RECT 0.6400 0.8000 1.6000 0.9000 ;
        RECT 1.5000 0.5150 1.6000 0.8000 ;
        RECT 0.6400 0.4700 0.7400 0.8000 ;
    END
    ANTENNADIFFAREA 0.266 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.2000 1.8200 1.8600 1.9200 ;
      RECT 1.7600 1.5050 1.8600 1.8200 ;
      RECT 0.1200 1.5150 1.3000 1.6150 ;
      RECT 1.2000 1.6150 1.3000 1.8200 ;
      RECT 0.1200 1.6150 0.2200 1.9450 ;
      RECT 0.6400 1.6150 0.7400 1.9450 ;
  END
END AOI21_X1P4M_A12TH

MACRO AOI21_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.6900 ;
        RECT 1.2000 0.3200 1.3000 0.6050 ;
        RECT 1.7600 0.3200 1.8600 0.6050 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4800 1.0500 1.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1542 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8300 1.3500 1.2500 ;
        RECT 1.2500 1.2500 1.6000 1.3500 ;
        RECT 0.6400 0.7300 1.6000 0.8300 ;
        RECT 1.5000 1.3500 1.6000 1.7000 ;
        RECT 1.5000 0.4250 1.6000 0.7300 ;
        RECT 0.6400 0.4200 0.7400 0.7300 ;
    END
    ANTENNADIFFAREA 0.375 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9300 0.3500 1.2500 ;
        RECT 0.2400 1.2500 1.1050 1.3500 ;
        RECT 1.0050 0.9500 1.1050 1.2500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.3800 1.7700 0.4800 2.0800 ;
        RECT 0.9000 1.7700 1.0000 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5050 1.0400 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.18 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 1.2000 1.8200 1.8600 1.9200 ;
      RECT 1.7600 1.5100 1.8600 1.8200 ;
      RECT 0.1200 1.5150 1.3000 1.6150 ;
      RECT 1.2000 1.6150 1.3000 1.8200 ;
      RECT 0.1200 1.6150 0.2200 1.9450 ;
      RECT 0.6400 1.6150 0.7400 1.9450 ;
  END
END AOI21_X2M_A12TH

MACRO AOI21_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6300 ;
        RECT 1.0800 0.3200 1.2500 0.5250 ;
        RECT 1.9350 0.3200 2.1050 0.5500 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 0.8500 1.5850 0.9400 ;
        RECT 0.4650 0.9400 1.5850 0.9500 ;
        RECT 0.4650 0.9500 0.8350 1.0400 ;
        RECT 1.4950 0.9500 1.5850 1.1000 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0100 1.0500 1.3800 1.1600 ;
        RECT 1.0100 1.1600 1.1000 1.2500 ;
        RECT 0.2350 1.2500 1.1000 1.3500 ;
        RECT 0.2350 1.0000 0.3250 1.2500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9000 1.0500 2.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 0.6500 2.3650 0.7500 ;
        RECT 1.7100 0.7500 1.8100 1.2600 ;
        RECT 0.5600 0.4600 0.7300 0.6500 ;
        RECT 2.1950 0.4600 2.3650 0.6500 ;
        RECT 1.6400 0.4500 1.8100 0.6500 ;
        RECT 1.7100 1.2600 2.5200 1.3500 ;
        RECT 1.9100 1.3500 2.0000 1.7000 ;
        RECT 2.4300 1.3500 2.5200 1.7200 ;
    END
    ANTENNADIFFAREA 0.70115 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.3400 1.7700 0.4300 2.0800 ;
        RECT 0.8600 1.7700 0.9500 2.0800 ;
        RECT 1.3900 1.7700 1.4800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6500 1.8300 2.2600 1.9200 ;
      RECT 2.1700 1.5000 2.2600 1.8300 ;
      RECT 0.0800 1.5300 1.7400 1.6300 ;
      RECT 1.6500 1.6300 1.7400 1.8300 ;
      RECT 0.0800 1.6400 0.1700 1.9600 ;
      RECT 0.6000 1.6400 0.6900 1.9600 ;
      RECT 0.0800 1.6300 1.2100 1.6400 ;
      RECT 1.1200 1.6400 1.2100 1.9600 ;
  END
END AOI21_X3M_A12TH

MACRO AOI21_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0550 0.3200 0.2250 0.5500 ;
        RECT 1.0950 0.3200 1.2650 0.5600 ;
        RECT 2.1500 0.3200 2.3200 0.5600 ;
        RECT 2.7100 0.3200 2.8000 0.5600 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7500 0.8500 1.5600 0.9500 ;
        RECT 1.4700 0.9500 1.5600 0.9700 ;
        RECT 0.7500 0.9500 0.8500 0.9600 ;
        RECT 1.4700 0.9700 1.8800 1.0600 ;
        RECT 0.4800 0.9600 0.8500 1.0600 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0000 1.0500 1.3800 1.1600 ;
        RECT 1.0000 1.1600 1.1000 1.2500 ;
        RECT 1.2900 1.1600 1.3800 1.2500 ;
        RECT 0.2500 1.2500 1.1000 1.3500 ;
        RECT 1.2900 1.2500 2.1250 1.3500 ;
        RECT 0.2500 1.0000 0.3400 1.2500 ;
        RECT 2.0350 1.0000 2.1250 1.2500 ;
    END
    ANTENNAGATEAREA 0.36 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5000 1.0500 2.9600 1.1500 ;
    END
    ANTENNAGATEAREA 0.3084 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5750 0.6500 2.5400 0.7500 ;
        RECT 2.2500 0.7500 2.5400 0.7800 ;
        RECT 1.6550 0.7500 1.7450 0.7800 ;
        RECT 0.5750 0.4600 0.7450 0.6500 ;
        RECT 1.6550 0.4100 1.7450 0.6500 ;
        RECT 2.4500 0.4100 2.5400 0.6500 ;
        RECT 2.2500 0.7800 2.3500 1.2500 ;
        RECT 2.2500 1.2500 3.0600 1.3500 ;
        RECT 2.4500 1.3500 2.5400 1.6350 ;
        RECT 2.9700 1.3500 3.0600 1.6350 ;
    END
    ANTENNADIFFAREA 0.75 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.3550 1.7700 0.4450 2.0800 ;
        RECT 0.8750 1.7700 0.9650 2.0800 ;
        RECT 1.3950 1.7700 1.4850 2.0800 ;
        RECT 1.9300 1.7700 2.0200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1900 1.8300 3.3200 1.9200 ;
      RECT 3.2300 1.5100 3.3200 1.8300 ;
      RECT 0.0950 1.5500 2.2800 1.6400 ;
      RECT 2.1900 1.6400 2.2800 1.8300 ;
      RECT 2.7100 1.5100 2.8000 1.8300 ;
      RECT 0.0950 1.6400 0.1850 1.9800 ;
      RECT 0.6150 1.6400 0.7050 1.9800 ;
      RECT 1.1350 1.6400 1.2250 1.9800 ;
      RECT 1.6550 1.6400 1.7450 1.9800 ;
  END
END AOI21_X4M_A12TH

MACRO AOI21_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.3800 0.3200 0.4800 0.7000 ;
        RECT 0.9000 0.3200 1.0000 0.7000 ;
        RECT 1.4200 0.3200 1.5200 0.7000 ;
        RECT 3.5900 0.3200 3.6900 0.6950 ;
        RECT 4.1100 0.3200 4.2100 0.6950 ;
        RECT 4.6400 0.3200 4.7400 0.6950 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9050 1.0350 3.1150 1.1500 ;
    END
    ANTENNAGATEAREA 0.54 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4700 1.0350 4.4800 1.1500 ;
    END
    ANTENNAGATEAREA 0.4632 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 0.9000 4.7500 1.3000 ;
        RECT 3.5000 1.3000 4.7500 1.4000 ;
        RECT 3.2550 0.8250 4.7500 0.9000 ;
        RECT 3.5000 1.4000 3.6000 1.7000 ;
        RECT 4.0200 1.4000 4.1200 1.7000 ;
        RECT 4.5400 1.4000 4.6400 1.7000 ;
        RECT 1.8850 0.8000 4.7500 0.8250 ;
        RECT 1.8850 0.7250 3.3550 0.8000 ;
        RECT 3.8500 0.4700 3.9500 0.8000 ;
        RECT 4.3800 0.4700 4.4800 0.8000 ;
    END
    ANTENNADIFFAREA 1.126 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3450 1.0350 1.5550 1.1500 ;
    END
    ANTENNAGATEAREA 0.54 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.3800 1.7700 0.4800 2.0800 ;
        RECT 0.9000 1.7700 1.0000 2.0800 ;
        RECT 1.4200 1.7700 1.5200 2.0800 ;
        RECT 1.9400 1.7700 2.0400 2.0800 ;
        RECT 2.4600 1.7700 2.5600 2.0800 ;
        RECT 2.9800 1.7700 3.0800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6800 0.4800 3.3950 0.5800 ;
      RECT 0.1200 0.8000 1.7800 0.9000 ;
      RECT 1.6800 0.5800 1.7800 0.8000 ;
      RECT 0.1200 0.4700 0.2200 0.8000 ;
      RECT 0.6400 0.4700 0.7400 0.8000 ;
      RECT 1.1600 0.4700 1.2600 0.8000 ;
      RECT 3.2400 1.8200 4.9000 1.9200 ;
      RECT 4.8000 1.5100 4.9000 1.8200 ;
      RECT 3.2400 1.4000 3.3400 1.8200 ;
      RECT 0.1200 1.3000 3.3400 1.4000 ;
      RECT 3.7600 1.5100 3.8600 1.8200 ;
      RECT 4.2800 1.5100 4.3800 1.8200 ;
      RECT 0.1200 1.4000 0.2200 1.7200 ;
      RECT 0.6400 1.4000 0.7400 1.7200 ;
      RECT 1.1600 1.4000 1.2600 1.7200 ;
      RECT 1.6800 1.4000 1.7800 1.7200 ;
      RECT 2.2000 1.4000 2.3000 1.7200 ;
      RECT 2.7200 1.4000 2.8200 1.7200 ;
  END
END AOI21_X6M_A12TH

MACRO AOI21_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.3800 0.3200 0.4800 0.6800 ;
        RECT 0.9000 0.3200 1.0000 0.6800 ;
        RECT 1.4200 0.3200 1.5200 0.6800 ;
        RECT 1.9400 0.3200 2.0400 0.6800 ;
        RECT 4.6300 0.3200 4.7300 0.6950 ;
        RECT 5.1750 0.3200 5.2750 0.6950 ;
        RECT 5.7250 0.3200 5.8250 0.6950 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3550 1.0350 2.0650 1.1500 ;
    END
    ANTENNAGATEAREA 0.72 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.3800 1.7900 0.4800 2.0800 ;
        RECT 0.9000 1.7900 1.0000 2.0800 ;
        RECT 1.4200 1.7900 1.5200 2.0800 ;
        RECT 1.9400 1.7900 2.0400 2.0800 ;
        RECT 2.4600 1.7900 2.5600 2.0800 ;
        RECT 2.9800 1.7900 3.0800 2.0800 ;
        RECT 3.5000 1.7900 3.6000 2.0800 ;
        RECT 4.0200 1.7900 4.1200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2350 0.9150 6.3650 1.2850 ;
        RECT 4.5250 1.2850 6.3650 1.4150 ;
        RECT 4.3200 0.8400 6.3650 0.9150 ;
        RECT 4.5250 1.4150 4.6550 1.7000 ;
        RECT 5.0450 1.4150 5.1750 1.7000 ;
        RECT 5.5650 1.4150 5.6950 1.7000 ;
        RECT 6.0850 1.4150 6.2150 1.7000 ;
        RECT 2.4050 0.7850 6.3650 0.8400 ;
        RECT 2.4050 0.7100 4.4500 0.7850 ;
        RECT 4.8750 0.4700 5.0050 0.7850 ;
        RECT 5.4450 0.4700 5.5750 0.7850 ;
        RECT 5.9750 0.4700 6.1050 0.7850 ;
    END
    ANTENNADIFFAREA 1.563 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5150 1.0350 6.0750 1.1500 ;
    END
    ANTENNAGATEAREA 0.6168 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4450 1.0350 4.1450 1.1500 ;
    END
    ANTENNAGATEAREA 0.72 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 2.2000 0.4800 4.4350 0.5800 ;
      RECT 0.1200 0.7800 2.3000 0.8800 ;
      RECT 2.2000 0.5800 2.3000 0.7800 ;
      RECT 0.1200 0.4700 0.2200 0.7800 ;
      RECT 0.6400 0.4700 0.7400 0.7800 ;
      RECT 1.1600 0.4700 1.2600 0.7800 ;
      RECT 1.6800 0.4700 1.7800 0.7800 ;
      RECT 4.2800 1.8200 6.4600 1.9200 ;
      RECT 6.3600 1.5200 6.4600 1.8200 ;
      RECT 4.2800 1.4000 4.3800 1.8200 ;
      RECT 0.1200 1.3000 4.3800 1.4000 ;
      RECT 4.8000 1.5100 4.9000 1.8200 ;
      RECT 5.3200 1.5100 5.4200 1.8200 ;
      RECT 5.8400 1.5100 5.9400 1.8200 ;
      RECT 0.1200 1.4000 0.2200 1.7150 ;
      RECT 0.6400 1.4000 0.7400 1.7000 ;
      RECT 1.1600 1.4000 1.2600 1.7000 ;
      RECT 1.6800 1.4000 1.7800 1.7000 ;
      RECT 2.2000 1.4000 2.3000 1.7000 ;
      RECT 2.7200 1.4000 2.8200 1.7000 ;
      RECT 3.2400 1.4000 3.3400 1.7000 ;
      RECT 3.7600 1.4000 3.8600 1.7000 ;
  END
END AOI21_X8M_A12TH

MACRO AOI221_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7200 ;
        RECT 1.0600 0.3200 1.1600 0.7100 ;
        RECT 1.6250 0.3200 1.7250 0.7200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.6900 0.9500 0.8000 ;
        RECT 0.8500 0.8000 1.5400 0.9000 ;
        RECT 0.5550 0.5900 0.9500 0.6900 ;
        RECT 1.4400 0.9000 1.5400 1.5450 ;
        RECT 1.3650 0.5200 1.4650 0.8000 ;
        RECT 1.3650 1.5450 1.5400 1.7150 ;
    END
    ANTENNADIFFAREA 0.1358 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6400 1.0350 1.7500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0363 ;
  END C0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8950 1.2500 1.3150 1.3500 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0250 0.5500 1.4350 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4350 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.3350 1.7850 0.4350 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.7500 1.0500 ;
        RECT 0.6500 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5700 1.2550 1.6700 ;
      RECT 0.5950 1.6700 0.6950 1.9900 ;
      RECT 0.0750 1.6700 0.1750 1.9900 ;
      RECT 0.8100 1.8200 1.7300 1.9200 ;
      RECT 1.6300 1.5300 1.7300 1.8200 ;
  END
END AOI221_X0P5M_A12TH

MACRO AOI221_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7100 ;
        RECT 1.0600 0.3200 1.1600 0.7050 ;
        RECT 1.6250 0.3200 1.7250 0.7100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.6950 0.9500 0.8000 ;
        RECT 0.8500 0.8000 1.5400 0.9000 ;
        RECT 0.5600 0.5950 0.9500 0.6950 ;
        RECT 1.4400 0.9000 1.5400 1.4750 ;
        RECT 1.3650 0.4900 1.4650 0.8000 ;
        RECT 1.3700 1.4750 1.5400 1.6450 ;
    END
    ANTENNADIFFAREA 0.1862 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.8100 0.7500 1.0500 ;
        RECT 0.6500 1.0500 0.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0400 0.5500 1.4600 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6400 1.0350 1.7500 1.4200 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END C0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4600 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.3000 1.7950 0.4700 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 1.2500 1.3200 1.3500 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END B1
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5850 1.2500 1.6850 ;
      RECT 0.5950 1.6850 0.6950 1.9900 ;
      RECT 0.0750 1.6850 0.1750 1.9900 ;
      RECT 0.8100 1.8200 1.7300 1.9200 ;
      RECT 1.6300 1.5300 1.7300 1.8200 ;
  END
END AOI221_X0P7M_A12TH

MACRO AOI221_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7200 ;
        RECT 1.0600 0.3200 1.1600 0.5300 ;
        RECT 1.6300 0.3200 1.7300 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.3350 1.7900 0.4350 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0400 0.5500 1.4750 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9000 0.8500 1.3200 0.9500 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4450 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6400 0.8550 1.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6650 1.0500 1.1600 1.1500 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 0.4100 0.7500 0.6200 ;
        RECT 0.5600 0.6200 1.5400 0.7200 ;
        RECT 1.4400 0.7200 1.5400 1.3000 ;
        RECT 1.3650 0.5150 1.4650 0.6200 ;
        RECT 1.3700 1.3000 1.5400 1.6700 ;
    END
    ANTENNADIFFAREA 0.2636 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5850 1.2150 1.6850 ;
      RECT 0.5950 1.6850 0.6950 1.9900 ;
      RECT 1.1150 1.3150 1.2150 1.5850 ;
      RECT 0.0750 1.6850 0.1750 1.9900 ;
      RECT 0.8100 1.8200 1.7300 1.9200 ;
      RECT 1.6300 1.5300 1.7300 1.8200 ;
  END
END AOI221_X1M_A12TH

MACRO AOI221_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0850 0.3200 0.1850 0.7050 ;
        RECT 1.1300 0.3200 1.2300 0.7050 ;
        RECT 1.4200 0.3200 1.5200 0.7050 ;
        RECT 2.4600 0.3200 2.5600 0.7050 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1150 1.2500 1.2050 1.3500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.2500 2.4500 1.3500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0500 0.8700 1.1500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5350 1.0500 2.9550 1.1500 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7950 1.0500 2.2150 1.1500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9000 3.1500 1.4500 ;
        RECT 2.7200 1.4500 3.1500 1.5500 ;
        RECT 0.6100 0.8000 3.1500 0.9000 ;
        RECT 2.7200 1.5500 2.8200 1.6900 ;
        RECT 2.7200 0.6350 2.8200 0.8000 ;
        RECT 0.6100 0.5700 0.7100 0.8000 ;
        RECT 1.9400 0.5700 2.0400 0.8000 ;
    END
    ANTENNADIFFAREA 0.31075 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.0900 1.6900 0.1900 2.0800 ;
        RECT 0.6100 1.6900 0.7100 2.0800 ;
        RECT 1.1300 1.6900 1.2300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3500 1.4400 2.3000 1.5400 ;
      RECT 1.6800 1.5400 1.7800 1.6650 ;
      RECT 2.2000 1.5400 2.3000 1.6650 ;
      RECT 0.3500 1.5400 0.4500 1.8850 ;
      RECT 0.8700 1.5400 0.9700 1.8850 ;
      RECT 1.3850 1.8200 3.1350 1.9200 ;
      RECT 1.3850 1.9200 1.5550 1.9250 ;
      RECT 1.9050 1.9200 2.0750 1.9250 ;
      RECT 2.4650 1.9200 2.5550 1.9250 ;
      RECT 1.3850 1.6350 1.5550 1.8200 ;
      RECT 1.9050 1.6350 2.0750 1.8200 ;
      RECT 2.4650 1.5350 2.5550 1.8200 ;
  END
END AOI221_X1P4M_A12TH

MACRO AOI221_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.6400 0.3200 0.7400 0.5700 ;
        RECT 1.6800 0.3200 1.7800 0.5700 ;
        RECT 2.4900 0.3200 2.5900 0.5600 ;
        RECT 3.0100 0.3200 3.1100 0.5700 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.2500 1.1050 1.3500 ;
        RECT 0.2000 1.1750 0.3000 1.2500 ;
        RECT 1.0050 1.0400 1.1050 1.2500 ;
        RECT 0.1300 1.0850 0.3000 1.1750 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3800 1.7900 0.4800 2.0800 ;
        RECT 0.9000 1.7900 1.0000 2.0800 ;
    END
  END VDD

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5400 1.0500 2.9600 1.1500 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0850 0.6600 2.8500 0.7600 ;
        RECT 2.2500 0.7600 2.3500 1.3000 ;
        RECT 2.7500 0.4400 2.8500 0.6600 ;
        RECT 0.0850 0.4200 0.2550 0.6600 ;
        RECT 1.1250 0.4200 1.2950 0.6600 ;
        RECT 2.1650 0.4200 2.3500 0.6600 ;
        RECT 2.2500 1.3000 2.8500 1.4000 ;
        RECT 2.7500 1.4000 2.8500 1.7000 ;
    END
    ANTENNADIFFAREA 0.4582 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 1.0400 2.1500 1.3000 ;
        RECT 1.2500 1.3000 2.1500 1.4000 ;
        RECT 1.2500 1.0400 1.3650 1.3000 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4900 1.0400 0.8900 1.1500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5300 1.0400 1.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END B1
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5100 2.3550 1.6100 ;
      RECT 1.1600 1.6100 1.2600 1.9400 ;
      RECT 0.1200 1.6100 0.2200 1.9400 ;
      RECT 0.6400 1.6100 0.7400 1.9400 ;
      RECT 1.3650 1.8200 3.1100 1.9200 ;
      RECT 3.0100 1.4900 3.1100 1.8200 ;
      RECT 2.4900 1.5100 2.5900 1.8200 ;
  END
END AOI221_X2M_A12TH

MACRO AOI221_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6100 ;
        RECT 1.1150 0.3200 1.2150 0.5600 ;
        RECT 2.1550 0.3200 2.2550 0.5600 ;
        RECT 3.1950 0.3200 3.2950 0.5600 ;
        RECT 3.4450 0.3200 3.5450 0.5600 ;
        RECT 3.9650 0.3200 4.0650 0.5600 ;
        RECT 0.0800 0.6100 0.1700 0.7600 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7400 1.3000 2.7500 1.4000 ;
        RECT 2.6400 1.1800 2.7500 1.3000 ;
        RECT 1.7400 1.0400 1.8400 1.3000 ;
        RECT 2.6400 1.0900 2.8300 1.1800 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 0.8350 1.1500 ;
        RECT 0.7350 0.9500 0.8350 1.0500 ;
        RECT 0.7350 0.8500 1.5800 0.9500 ;
        RECT 1.4800 0.9500 1.5800 1.1550 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.6950 1.0500 4.1200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END C0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1500 1.2500 1.1550 1.3500 ;
        RECT 0.1500 1.1850 0.2500 1.2500 ;
        RECT 1.0550 1.1800 1.1550 1.2500 ;
        RECT 0.0500 1.0850 0.2500 1.1850 ;
        RECT 1.0550 1.0900 1.2700 1.1800 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.7500 3.5500 1.2900 ;
        RECT 3.4500 1.2900 4.3250 1.3900 ;
        RECT 0.5600 0.6500 4.3250 0.7500 ;
        RECT 3.7050 1.3900 3.8050 1.7000 ;
        RECT 4.2250 1.3900 4.3250 1.7200 ;
        RECT 3.7050 0.4400 3.8050 0.6500 ;
        RECT 4.2250 0.4400 4.3250 0.6500 ;
        RECT 0.5600 0.4100 0.7300 0.6500 ;
        RECT 1.6000 0.4100 1.7700 0.6500 ;
        RECT 2.6400 0.4100 2.8100 0.6500 ;
    END
    ANTENNADIFFAREA 0.6516 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 0.3350 1.7700 0.4350 2.0800 ;
        RECT 0.8550 1.7700 0.9550 2.0800 ;
        RECT 1.3750 1.7700 1.4750 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0200 1.0500 2.3950 1.1500 ;
        RECT 2.2950 0.9500 2.3950 1.0500 ;
        RECT 2.2950 0.8500 3.1150 0.9500 ;
        RECT 3.0150 0.9500 3.1150 1.1450 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B1
  OBS
    LAYER M1 ;
      RECT 0.0750 1.5100 3.3500 1.6100 ;
      RECT 1.6350 1.6100 1.7350 1.9400 ;
      RECT 0.0750 1.6100 0.1750 1.9400 ;
      RECT 0.5950 1.6100 0.6950 1.9400 ;
      RECT 1.1150 1.6100 1.2150 1.9400 ;
      RECT 1.8450 1.8200 4.0650 1.9200 ;
      RECT 3.9650 1.5100 4.0650 1.8200 ;
      RECT 3.4450 1.5100 3.5450 1.8200 ;
  END
END AOI221_X3M_A12TH

MACRO AOI221_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.6100 0.3200 0.7100 0.5600 ;
        RECT 1.6500 0.3200 1.7500 0.5600 ;
        RECT 2.6900 0.3200 2.7900 0.5600 ;
        RECT 3.7300 0.3200 3.8300 0.5600 ;
        RECT 4.5400 0.3200 4.6400 0.5600 ;
        RECT 5.0600 0.3200 5.1600 0.5600 ;
        RECT 5.5800 0.3200 5.6800 0.6100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7500 4.5500 1.2900 ;
        RECT 4.4500 1.2900 5.4200 1.3900 ;
        RECT 0.0550 0.6500 5.4200 0.7500 ;
        RECT 4.8000 1.3900 4.9000 1.7000 ;
        RECT 5.3200 1.3900 5.4200 1.7000 ;
        RECT 4.8000 0.4400 4.9000 0.6500 ;
        RECT 5.3200 0.4400 5.4200 0.6500 ;
        RECT 0.0550 0.4100 0.2250 0.6500 ;
        RECT 1.0950 0.4100 1.2650 0.6500 ;
        RECT 2.1350 0.4100 2.3050 0.6500 ;
        RECT 3.1750 0.4100 3.3450 0.6500 ;
        RECT 4.2150 0.4100 4.3850 0.6500 ;
    END
    ANTENNADIFFAREA 0.8345 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4750 1.0500 0.8500 1.1500 ;
        RECT 0.7500 0.9500 0.8500 1.0500 ;
        RECT 0.7500 0.8500 1.6100 0.9500 ;
        RECT 1.5100 0.9500 1.6100 1.0500 ;
        RECT 1.5100 1.0500 1.8850 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8400 1.0500 5.3600 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END C0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 1.3900 1.7700 1.4900 2.0800 ;
        RECT 1.9100 1.7700 2.0100 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2000 1.2900 2.1150 1.3900 ;
        RECT 0.2000 1.1450 0.3000 1.2900 ;
        RECT 1.0500 1.0900 1.2850 1.2900 ;
        RECT 2.0150 1.0400 2.1150 1.2900 ;
        RECT 0.1250 1.0450 0.3000 1.1450 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5500 1.0500 2.9300 1.1500 ;
        RECT 2.8300 0.9500 2.9300 1.0500 ;
        RECT 2.8300 0.8500 3.6900 0.9500 ;
        RECT 3.5900 0.9500 3.6900 1.0500 ;
        RECT 3.5900 1.0500 3.9650 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2800 1.2950 4.1900 1.3850 ;
        RECT 4.1000 1.1700 4.1900 1.2950 ;
        RECT 3.1550 1.0900 3.3900 1.2950 ;
        RECT 2.2800 1.0400 2.3700 1.2950 ;
        RECT 4.1000 1.0800 4.2800 1.1700 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.0900 1.5050 4.4050 1.6050 ;
      RECT 2.1700 1.6050 2.2700 1.9350 ;
      RECT 0.0900 1.6050 0.1900 1.9350 ;
      RECT 0.6100 1.6050 0.7100 1.9350 ;
      RECT 1.1300 1.6050 1.2300 1.9350 ;
      RECT 1.6500 1.6050 1.7500 1.9350 ;
      RECT 2.3750 1.8200 5.6800 1.9200 ;
      RECT 5.5800 1.4900 5.6800 1.8200 ;
      RECT 4.5400 1.5100 4.6400 1.8200 ;
      RECT 5.0600 1.5100 5.1600 1.8200 ;
  END
END AOI221_X4M_A12TH

MACRO AOI222_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7150 ;
        RECT 1.1350 0.3200 1.2350 0.7150 ;
        RECT 1.9700 0.3200 2.0700 0.7200 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0000 0.9100 1.1000 ;
        RECT 0.6500 1.1000 0.7500 1.3050 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0000 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.0000 1.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END B1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.0000 1.5550 1.4000 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END C0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9650 1.9600 1.3900 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.8100 1.7500 0.9100 ;
        RECT 1.6500 0.9100 1.7500 1.4900 ;
        RECT 0.6150 0.5550 0.7150 0.8100 ;
        RECT 1.4350 0.5400 1.5350 0.8100 ;
        RECT 1.6500 1.4900 1.8250 1.6600 ;
    END
    ANTENNADIFFAREA 0.171925 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.3550 1.7050 0.4550 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5150 1.2900 1.6050 ;
      RECT 0.6150 1.6050 0.7150 1.9300 ;
      RECT 0.0950 1.6050 0.1950 1.9300 ;
      RECT 0.8400 1.8100 2.0700 1.9000 ;
      RECT 1.9700 1.4900 2.0700 1.8100 ;
      RECT 1.4350 1.4900 1.5350 1.8100 ;
  END
END AOI222_X0P5M_A12TH

MACRO AOI222_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7200 ;
        RECT 1.1350 0.3200 1.2350 0.7200 ;
        RECT 1.9700 0.3200 2.0700 0.7200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.3550 1.7050 0.4550 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0000 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.0000 1.5550 1.4000 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END C0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.0000 1.1500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0000 0.9050 1.1000 ;
        RECT 0.6500 1.1000 0.7500 1.3050 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END B0

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.9650 1.9600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.8100 1.7500 0.9100 ;
        RECT 1.6500 0.9100 1.7500 1.4900 ;
        RECT 0.6150 0.5900 0.7150 0.8100 ;
        RECT 1.4350 0.5750 1.5350 0.8100 ;
        RECT 1.6500 1.4900 1.8250 1.6600 ;
    END
    ANTENNADIFFAREA 0.243175 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5150 1.2900 1.6050 ;
      RECT 0.6150 1.6050 0.7150 1.9450 ;
      RECT 0.0950 1.6050 0.1950 1.9450 ;
      RECT 0.8400 1.8300 2.0700 1.9200 ;
      RECT 1.9700 1.5100 2.0700 1.8300 ;
      RECT 1.4350 1.5100 1.5350 1.8300 ;
  END
END AOI222_X0P7M_A12TH

MACRO AOI222_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.7200 ;
        RECT 1.1350 0.3200 1.2350 0.7200 ;
        RECT 1.9700 0.3200 2.0700 0.7200 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.8950 0.1600 1.3050 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0000 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6150 0.8100 1.7500 0.9100 ;
        RECT 1.6500 0.9100 1.7500 1.3700 ;
        RECT 0.6150 0.4100 0.7150 0.8100 ;
        RECT 1.4350 0.4100 1.5350 0.8100 ;
        RECT 1.6500 1.3700 1.7950 1.7400 ;
    END
    ANTENNADIFFAREA 0.34385 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.0000 1.5550 1.4000 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END C0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.3550 1.7900 0.4550 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0000 0.9050 1.1000 ;
        RECT 0.6500 1.1000 0.7500 1.3050 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 1.0000 1.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8100 1.9600 1.2600 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END C1
  OBS
    LAYER M1 ;
      RECT 0.0950 1.4800 1.2900 1.5700 ;
      RECT 0.6150 1.5700 0.7150 1.9100 ;
      RECT 0.0950 1.5700 0.1950 1.9100 ;
      RECT 0.8200 1.8300 2.0700 1.9200 ;
      RECT 1.9700 1.4900 2.0700 1.8300 ;
      RECT 1.4350 1.5000 1.5350 1.8300 ;
  END
END AOI222_X1M_A12TH

MACRO AOI222_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.1600 0.3200 0.2500 0.5800 ;
        RECT 1.8300 0.3200 2.0000 0.5050 ;
        RECT 2.3550 0.3200 2.5250 0.5050 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.6850 1.4800 0.7500 ;
        RECT 0.6600 0.6500 3.0450 0.6850 ;
        RECT 2.3300 0.6850 2.4200 1.4400 ;
        RECT 2.8750 0.6850 3.0450 0.7000 ;
        RECT 0.6600 0.4500 0.8300 0.6500 ;
        RECT 1.3100 0.5950 3.0450 0.6500 ;
        RECT 2.3300 1.4400 3.3000 1.5300 ;
        RECT 1.3100 0.4300 1.4800 0.5950 ;
        RECT 2.8750 0.4100 3.0450 0.5950 ;
        RECT 2.6100 1.5300 2.7800 1.7300 ;
        RECT 3.1300 1.5300 3.3000 1.7300 ;
    END
    ANTENNADIFFAREA 0.59625 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7450 1.0500 3.1200 1.1700 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END C0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.8100 1.7500 0.9950 ;
        RECT 1.6500 0.9950 1.9400 1.0950 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2650 0.8500 1.1900 0.9500 ;
        RECT 0.2650 0.9500 0.3550 1.0700 ;
        RECT 1.1000 0.9500 1.1900 1.0800 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5100 1.2600 3.4100 1.3500 ;
        RECT 3.2100 1.2500 3.4100 1.2600 ;
        RECT 2.5100 0.9400 2.6000 1.2600 ;
        RECT 3.3200 1.2100 3.4100 1.2500 ;
        RECT 2.5100 0.8500 2.7000 0.9400 ;
        RECT 3.3200 1.1200 3.5250 1.2100 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END C1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.8750 2.1500 1.1850 ;
        RECT 1.4500 1.1850 2.1500 1.2750 ;
        RECT 2.0500 0.7750 2.2200 0.8750 ;
        RECT 1.4500 1.0400 1.5500 1.1850 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0500 0.9900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 1.1300 1.9500 1.2200 2.0800 ;
        RECT 0.0800 1.8200 0.1700 2.0800 ;
        RECT 0.6000 1.8200 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 1.4550 1.2000 1.5500 ;
      RECT 0.8600 1.5500 0.9500 1.9450 ;
      RECT 0.3400 1.4500 2.2200 1.4550 ;
      RECT 1.6100 1.4550 1.7000 1.7350 ;
      RECT 2.1300 1.4550 2.2200 1.7350 ;
      RECT 1.1000 1.3650 2.2200 1.4500 ;
      RECT 0.3400 1.5500 0.4300 1.9450 ;
      RECT 1.4000 1.8350 3.5200 1.9150 ;
      RECT 1.3100 1.8250 3.5200 1.8350 ;
      RECT 3.4300 1.5450 3.5200 1.8250 ;
      RECT 2.3900 1.9150 2.4800 1.9900 ;
      RECT 2.3900 1.6200 2.4800 1.8250 ;
      RECT 1.3100 1.5450 1.4900 1.8250 ;
      RECT 1.8700 1.5450 1.9600 1.8250 ;
      RECT 2.9100 1.9150 3.0000 1.9900 ;
      RECT 2.9100 1.6200 3.0000 1.8250 ;
  END
END AOI222_X1P4M_A12TH

MACRO AOI222_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.5750 0.3200 0.7450 0.5050 ;
        RECT 1.6150 0.3200 1.7850 0.5250 ;
        RECT 3.2300 0.3200 3.3300 0.6600 ;
    END
  END VSS

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1000 1.0500 3.6000 1.1600 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END C1

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 1.0350 2.9900 1.1650 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END C0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 1.0300 1.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END B1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9800 2.1600 1.2500 ;
        RECT 1.2350 1.2500 2.1600 1.3500 ;
        RECT 1.2350 0.9750 1.3350 1.2500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0250 0.8650 1.1550 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2500 1.0750 1.3500 ;
        RECT 0.2400 0.9950 0.3500 1.2500 ;
        RECT 0.9750 0.9750 1.0750 1.2500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7500 2.3500 1.3000 ;
        RECT 2.2500 1.3000 3.5900 1.4000 ;
        RECT 2.1000 0.7200 2.8450 0.7500 ;
        RECT 2.4550 1.4000 2.5450 1.6900 ;
        RECT 2.9700 1.4000 3.0700 1.7100 ;
        RECT 3.4900 1.4000 3.5900 1.7500 ;
        RECT 0.0550 0.6600 2.8450 0.7200 ;
        RECT 0.0550 0.6200 2.3050 0.6600 ;
        RECT 0.0550 0.4300 0.2250 0.6200 ;
        RECT 1.0950 0.4300 1.2650 0.6200 ;
    END
    ANTENNADIFFAREA 0.793 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0900 1.5500 2.3250 1.6400 ;
      RECT 1.1300 1.6400 1.2300 1.9800 ;
      RECT 0.0900 1.6400 0.1900 1.9800 ;
      RECT 0.6100 1.6400 0.7100 1.9800 ;
      RECT 1.3400 1.8300 3.3300 1.9200 ;
      RECT 3.2300 1.5100 3.3300 1.8300 ;
      RECT 2.7100 1.5100 2.8100 1.8300 ;
      RECT 2.9700 0.7600 3.5900 0.8500 ;
      RECT 3.4900 0.4500 3.5900 0.7600 ;
      RECT 2.9700 0.5700 3.0700 0.7600 ;
      RECT 2.4150 0.4800 3.0700 0.5700 ;
  END
END AOI222_X2M_A12TH

MACRO AO21_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 1.1750 0.3200 1.2650 0.4800 ;
        RECT 0.0950 0.3200 0.1850 0.8500 ;
        RECT 0.8550 0.4800 1.2650 0.5700 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3150 1.7200 0.4850 2.0800 ;
        RECT 1.1500 1.6000 1.2400 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 0.5400 1.5500 0.9700 ;
        RECT 1.4500 0.9700 1.5500 1.3850 ;
        RECT 1.4100 1.3850 1.5500 1.8150 ;
    END
    ANTENNADIFFAREA 0.202125 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1500 1.3900 ;
        RECT 0.0500 1.0000 0.2950 1.1000 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6900 1.0400 1.0400 1.1600 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9600 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5100 0.7050 1.6000 ;
      RECT 0.6150 1.6000 0.7050 1.9400 ;
      RECT 0.0950 1.6000 0.1850 1.9400 ;
      RECT 0.8800 1.4100 1.2700 1.5000 ;
      RECT 1.1800 0.7600 1.2700 1.4100 ;
      RECT 0.6150 0.6700 1.2700 0.7600 ;
      RECT 0.8800 1.5000 0.9700 1.8800 ;
      RECT 0.6150 0.4900 0.7050 0.6700 ;
  END
END AO21_X0P7M_A12TH

MACRO AO21_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.7600 ;
        RECT 0.8700 0.3200 0.9700 0.5700 ;
        RECT 1.1550 0.3200 1.2450 0.6400 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1450 1.7700 1.2350 2.0800 ;
        RECT 0.3550 1.7200 0.4450 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 0.5400 1.5500 0.9700 ;
        RECT 1.4500 0.9700 1.5500 1.2900 ;
        RECT 1.4100 1.2900 1.5500 1.7200 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1500 1.3900 ;
        RECT 0.0500 1.0000 0.2950 1.1000 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6700 1.0450 1.0650 1.1550 ;
    END
    ANTENNAGATEAREA 0.0633 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0050 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0738 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5100 0.7050 1.6000 ;
      RECT 0.6150 1.6000 0.7050 1.9400 ;
      RECT 0.0950 1.6000 0.1850 1.9400 ;
      RECT 0.8750 1.4800 1.2750 1.5700 ;
      RECT 1.1850 0.8500 1.2750 1.4800 ;
      RECT 0.5900 0.7600 1.2750 0.8500 ;
      RECT 0.5900 0.4600 0.6800 0.7600 ;
      RECT 0.8750 1.5700 0.9650 1.9100 ;
  END
END AO21_X1M_A12TH

MACRO AO21_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7600 ;
        RECT 1.0650 0.3200 1.2750 0.5100 ;
        RECT 1.7400 0.3200 1.9500 0.5100 ;
        RECT 2.4300 0.3200 2.5200 0.7600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.3400 1.6900 0.4300 2.0800 ;
        RECT 0.8600 1.6900 0.9500 2.0800 ;
        RECT 2.4300 1.6800 2.5200 2.0800 ;
        RECT 1.9100 1.6400 2.0000 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9500 2.5500 1.4500 ;
        RECT 2.1650 1.4500 2.5500 1.5500 ;
        RECT 2.1650 0.8500 2.5500 0.9500 ;
        RECT 2.1650 1.5500 2.2650 1.8800 ;
        RECT 2.1650 0.4800 2.2650 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0200 0.9500 1.1500 1.2350 ;
        RECT 0.1800 0.8500 1.1500 0.9500 ;
    END
    ANTENNAGATEAREA 0.1068 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2600 1.0500 1.6800 1.1500 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 0.8800 1.1500 ;
    END
    ANTENNAGATEAREA 0.1068 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0800 1.4800 1.2100 1.5700 ;
      RECT 1.1200 1.5700 1.2100 1.8300 ;
      RECT 1.1200 1.8300 1.7450 1.9200 ;
      RECT 1.6550 1.4900 1.7450 1.8300 ;
      RECT 0.0800 1.5700 0.1700 1.9000 ;
      RECT 0.6000 1.5700 0.6900 1.9000 ;
      RECT 1.8550 1.0700 2.3500 1.1600 ;
      RECT 1.3950 1.3000 1.9450 1.3900 ;
      RECT 1.8550 1.1600 1.9450 1.3000 ;
      RECT 1.8550 0.7200 1.9450 1.0700 ;
      RECT 0.6000 0.6300 1.9450 0.7200 ;
      RECT 0.6000 0.5100 0.6900 0.6300 ;
      RECT 1.3950 1.3900 1.4850 1.7100 ;
      RECT 1.3950 0.4400 1.4850 0.6300 ;
  END
END AO21_X1P4M_A12TH

MACRO AO21_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7600 ;
        RECT 1.1250 0.3200 1.2250 0.5350 ;
        RECT 1.6500 0.3200 1.7500 0.5350 ;
        RECT 1.9100 0.3200 2.0000 0.6850 ;
        RECT 2.4300 0.3200 2.5200 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 1.9100 1.7700 2.0000 2.0800 ;
        RECT 2.4300 1.7700 2.5200 2.0800 ;
        RECT 0.3400 1.6900 0.4300 2.0800 ;
        RECT 0.8600 1.6900 0.9500 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 0.9500 2.5500 1.2900 ;
        RECT 2.1650 1.2900 2.5500 1.3900 ;
        RECT 2.1650 0.8500 2.5500 0.9500 ;
        RECT 2.1650 1.3900 2.2650 1.7200 ;
        RECT 2.1650 0.5200 2.2650 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9500 0.3500 1.1900 ;
        RECT 0.2500 0.8500 1.0600 0.9500 ;
        RECT 0.9600 0.9500 1.0600 1.1900 ;
    END
    ANTENNAGATEAREA 0.1404 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1900 1.0500 1.6100 1.1500 ;
    END
    ANTENNAGATEAREA 0.12 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0450 0.8400 1.1550 ;
    END
    ANTENNAGATEAREA 0.1404 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0800 1.4800 1.2100 1.5700 ;
      RECT 1.1200 1.5700 1.2100 1.8300 ;
      RECT 1.1200 1.8300 1.7450 1.9200 ;
      RECT 1.6550 1.4900 1.7450 1.8300 ;
      RECT 0.0800 1.5700 0.1700 1.9100 ;
      RECT 0.6000 1.5700 0.6900 1.9100 ;
      RECT 1.7000 1.0800 2.3600 1.1700 ;
      RECT 0.5600 0.4550 0.7300 0.6550 ;
      RECT 1.3950 1.3900 1.4850 1.7100 ;
      RECT 1.3950 0.4400 1.4850 0.6550 ;
      RECT 1.3950 1.3000 1.7900 1.3900 ;
      RECT 1.7000 1.1700 1.7900 1.3000 ;
      RECT 1.7000 0.7450 1.7900 1.0800 ;
      RECT 0.5600 0.6550 1.7900 0.7450 ;
  END
END AO21_X2M_A12TH

MACRO AO21_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.8450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.6800 ;
        RECT 1.1250 0.3200 1.2950 0.5550 ;
        RECT 1.9000 0.3200 2.1100 0.5300 ;
        RECT 2.4200 0.3200 2.6300 0.5300 ;
        RECT 2.8050 0.3200 2.8950 0.6850 ;
        RECT 3.3250 0.3200 3.4150 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.8450 2.7200 ;
        RECT 2.8050 1.7700 2.8950 2.0800 ;
        RECT 3.3250 1.7700 3.4150 2.0800 ;
        RECT 0.3850 1.6900 0.4750 2.0800 ;
        RECT 0.9050 1.6900 0.9950 2.0800 ;
        RECT 1.4250 1.6900 1.5150 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0600 0.8500 3.6800 0.9500 ;
        RECT 3.4500 0.9500 3.5500 1.2900 ;
        RECT 3.0600 0.5200 3.1600 0.8500 ;
        RECT 3.5800 0.5200 3.6800 0.8500 ;
        RECT 3.0600 1.2900 3.6800 1.3900 ;
        RECT 3.0600 1.3900 3.1600 1.7200 ;
        RECT 3.5800 1.3900 3.6800 1.7200 ;
    END
    ANTENNADIFFAREA 0.658125 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2200 0.8500 1.4150 0.9500 ;
    END
    ANTENNAGATEAREA 0.2124 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8700 1.0500 2.3800 1.1500 ;
    END
    ANTENNAGATEAREA 0.1818 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 0.8800 1.7500 1.2500 ;
        RECT 0.8200 1.2500 1.7500 1.3500 ;
        RECT 0.8200 1.1500 0.9200 1.2500 ;
        RECT 0.5100 1.0500 0.9200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2124 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.1250 1.4800 1.7900 1.5700 ;
      RECT 1.6850 1.5700 1.7900 1.8300 ;
      RECT 1.6850 1.8300 2.3100 1.9200 ;
      RECT 2.2200 1.4900 2.3100 1.8300 ;
      RECT 0.1250 1.5700 0.2150 1.9100 ;
      RECT 0.6450 1.5700 0.7350 1.9100 ;
      RECT 1.1650 1.5700 1.2550 1.9100 ;
      RECT 2.5950 1.0800 3.3300 1.1700 ;
      RECT 0.6050 0.4100 0.7750 0.6500 ;
      RECT 1.6850 0.5050 1.7750 0.6500 ;
      RECT 1.9600 1.3900 2.0500 1.7100 ;
      RECT 2.2200 0.5050 2.3100 0.6500 ;
      RECT 1.9600 1.3000 2.6850 1.3900 ;
      RECT 2.4800 1.3900 2.5700 1.7800 ;
      RECT 2.5950 1.1700 2.6850 1.3000 ;
      RECT 2.5950 0.7400 2.6850 1.0800 ;
      RECT 0.6050 0.6500 2.6850 0.7400 ;
  END
END AO21_X3M_A12TH

MACRO AO21_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.0450 0.3200 ;
        RECT 0.1250 0.3200 0.2150 0.6300 ;
        RECT 1.1650 0.3200 1.2550 0.5800 ;
        RECT 1.9200 0.3200 2.0900 0.5350 ;
        RECT 2.4400 0.3200 2.6100 0.5350 ;
        RECT 2.7750 0.3200 2.8650 0.6850 ;
        RECT 3.2950 0.3200 3.3850 0.6850 ;
        RECT 3.8150 0.3200 3.9050 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.0450 2.7200 ;
        RECT 0.3850 1.7700 0.4750 2.0800 ;
        RECT 0.9050 1.7700 0.9950 2.0800 ;
        RECT 1.4250 1.7700 1.5150 2.0800 ;
        RECT 2.7750 1.7700 2.8650 2.0800 ;
        RECT 3.2950 1.7700 3.3850 2.0800 ;
        RECT 3.8150 1.7700 3.9050 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0300 0.8500 3.7500 0.9500 ;
        RECT 3.6500 0.9500 3.7500 1.3000 ;
        RECT 3.5550 0.5400 3.6450 0.8500 ;
        RECT 3.0300 0.5200 3.1300 0.8500 ;
        RECT 3.0300 1.3000 3.7500 1.4000 ;
        RECT 3.0300 1.4000 3.1300 1.7300 ;
        RECT 3.5550 1.4000 3.6450 1.7300 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 0.9500 0.3500 1.1900 ;
        RECT 0.2300 0.8500 1.1300 0.9500 ;
        RECT 1.0400 0.9500 1.4500 1.0400 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8700 1.0500 2.3900 1.1500 ;
    END
    ANTENNAGATEAREA 0.2313 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6200 0.9800 1.7500 1.2500 ;
        RECT 0.8200 1.2500 1.7500 1.3500 ;
        RECT 0.8200 1.1500 0.9200 1.2500 ;
        RECT 0.5100 1.0500 0.9200 1.1500 ;
    END
    ANTENNAGATEAREA 0.27 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.1250 1.4800 1.7750 1.5700 ;
      RECT 1.6850 1.5700 1.7750 1.8300 ;
      RECT 1.6850 1.8300 2.3100 1.9200 ;
      RECT 2.2200 1.4900 2.3100 1.8300 ;
      RECT 0.1250 1.5700 0.2150 1.9100 ;
      RECT 0.6450 1.5700 0.7350 1.9100 ;
      RECT 1.1650 1.5700 1.2550 1.9100 ;
      RECT 2.5650 1.0900 3.4800 1.1800 ;
      RECT 0.6050 0.4700 0.7750 0.6700 ;
      RECT 1.6450 0.4700 1.8150 0.6700 ;
      RECT 1.9600 1.3900 2.0500 1.7000 ;
      RECT 2.1800 0.4700 2.3500 0.6700 ;
      RECT 1.9600 1.3000 2.6550 1.3900 ;
      RECT 2.4800 1.3900 2.5700 1.7200 ;
      RECT 2.5650 1.1800 2.6550 1.3000 ;
      RECT 2.5650 0.7600 2.6550 1.0900 ;
      RECT 0.6050 0.6700 2.6550 0.7600 ;
  END
END AO21_X4M_A12TH

MACRO AO21_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1850 0.6700 ;
        RECT 1.0950 0.3200 1.2650 0.5450 ;
        RECT 2.1350 0.3200 2.3050 0.5450 ;
        RECT 2.9300 0.3200 3.1000 0.5550 ;
        RECT 3.4500 0.3200 3.6200 0.5550 ;
        RECT 3.9700 0.3200 4.1400 0.5550 ;
        RECT 4.2600 0.3200 4.3500 0.6850 ;
        RECT 4.7800 0.3200 4.8700 0.6850 ;
        RECT 5.3000 0.3200 5.3900 0.6850 ;
        RECT 5.8200 0.3200 5.9100 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 4.2600 1.7700 4.3500 2.0800 ;
        RECT 4.7800 1.7700 4.8700 2.0800 ;
        RECT 5.3000 1.7700 5.3900 2.0800 ;
        RECT 5.8200 1.7700 5.9100 2.0800 ;
        RECT 0.3550 1.7350 0.4450 2.0800 ;
        RECT 0.8750 1.7350 0.9650 2.0800 ;
        RECT 1.3950 1.7350 1.4850 2.0800 ;
        RECT 1.9150 1.7350 2.0050 2.0800 ;
        RECT 2.4350 1.7300 2.5250 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5150 0.8500 5.6500 0.9500 ;
        RECT 5.4500 0.9500 5.5500 1.2900 ;
        RECT 5.5600 0.5400 5.6500 0.8500 ;
        RECT 4.5150 0.5200 4.6150 0.8500 ;
        RECT 5.0400 0.5200 5.1300 0.8500 ;
        RECT 4.5150 1.2900 5.6500 1.3900 ;
        RECT 4.5150 1.3900 4.6150 1.7200 ;
        RECT 5.0400 1.3900 5.1300 1.7200 ;
        RECT 5.5600 1.3900 5.6500 1.7200 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9500 0.3500 1.1900 ;
        RECT 0.2500 0.8500 2.4000 0.9500 ;
        RECT 0.9900 0.9500 1.3600 1.0100 ;
        RECT 2.0300 0.9500 2.4000 1.0100 ;
    END
    ANTENNAGATEAREA 0.4155 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9500 1.0500 3.8650 1.1500 ;
    END
    ANTENNAGATEAREA 0.3555 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5900 1.0050 2.7500 1.2500 ;
        RECT 0.7700 1.2500 2.7500 1.3500 ;
        RECT 0.7700 1.1500 0.8700 1.2500 ;
        RECT 1.5200 1.0950 1.8900 1.2500 ;
        RECT 0.4700 1.0500 0.8700 1.1500 ;
    END
    ANTENNAGATEAREA 0.4155 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0950 1.4800 2.7850 1.5700 ;
      RECT 2.6950 1.5700 2.7850 1.8300 ;
      RECT 2.6950 1.8300 3.8400 1.9200 ;
      RECT 3.2300 1.4900 3.3200 1.8300 ;
      RECT 3.7500 1.4900 3.8400 1.8300 ;
      RECT 0.0950 1.5700 0.1850 1.9100 ;
      RECT 0.6150 1.5700 0.7050 1.9100 ;
      RECT 1.1350 1.5700 1.2250 1.9100 ;
      RECT 1.6550 1.5700 1.7450 1.9100 ;
      RECT 2.1750 1.5700 2.2650 1.9100 ;
      RECT 4.0100 1.0800 5.3250 1.1700 ;
      RECT 0.5750 0.4500 0.7450 0.6500 ;
      RECT 1.6150 0.4500 1.7850 0.6500 ;
      RECT 2.6550 0.4500 2.8250 0.6500 ;
      RECT 2.9700 1.3700 3.0600 1.7100 ;
      RECT 3.1900 0.4500 3.3600 0.6500 ;
      RECT 3.4900 1.3700 3.5800 1.7100 ;
      RECT 3.7100 0.4500 3.8800 0.6500 ;
      RECT 2.9700 1.2800 4.1000 1.3700 ;
      RECT 4.0100 1.3700 4.1000 1.7100 ;
      RECT 4.0100 1.1700 4.1000 1.2800 ;
      RECT 4.0100 0.7400 4.1000 1.0800 ;
      RECT 0.5750 0.6500 4.1000 0.7400 ;
  END
END AO21_X6M_A12TH

MACRO AO22_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7500 ;
        RECT 1.1150 0.3200 1.2150 0.7200 ;
        RECT 1.3700 0.3200 1.4600 0.9200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.3400 1.7600 0.4300 2.0800 ;
        RECT 1.3700 1.5200 1.4600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9200 1.7500 1.4950 ;
        RECT 1.6250 1.4950 1.7500 1.9250 ;
        RECT 1.6250 0.5100 1.7500 0.9200 ;
    END
    ANTENNADIFFAREA 0.1304 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0050 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8400 1.1700 1.1900 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0400 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END A0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 0.9350 0.7650 1.3350 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END B0
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5100 0.6900 1.6000 ;
      RECT 0.6000 1.6000 0.6900 1.8300 ;
      RECT 0.6000 1.8300 1.2100 1.9200 ;
      RECT 1.1200 1.5100 1.2100 1.8300 ;
      RECT 0.0800 1.6000 0.1700 1.9400 ;
      RECT 0.8600 1.3000 1.5400 1.3900 ;
      RECT 1.4500 1.0200 1.5400 1.3000 ;
      RECT 0.8600 1.3900 0.9500 1.7100 ;
      RECT 0.8600 0.7000 0.9500 1.3000 ;
      RECT 0.5400 0.6100 0.9500 0.7000 ;
  END
END AO22_X0P5M_A12TH

MACRO AO22_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.8800 ;
        RECT 1.1100 0.3200 1.2200 0.7050 ;
        RECT 1.3700 0.3200 1.4600 0.8700 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0000 0.1600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0400 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8300 1.1700 1.1900 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.3000 1.7200 0.4700 2.0800 ;
        RECT 1.3700 1.5950 1.4600 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0100 0.7650 1.3600 ;
    END
    ANTENNAGATEAREA 0.0585 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9200 1.7500 1.4900 ;
        RECT 1.6300 1.4900 1.7500 1.9200 ;
        RECT 1.6300 0.5100 1.7500 0.9200 ;
    END
    ANTENNADIFFAREA 0.1848 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5100 0.6900 1.6000 ;
      RECT 0.6000 1.6000 0.6900 1.8300 ;
      RECT 0.6000 1.8300 1.2100 1.9200 ;
      RECT 1.1200 1.5100 1.2100 1.8300 ;
      RECT 0.0800 1.6000 0.1700 1.9400 ;
      RECT 0.8600 1.3000 1.5500 1.3900 ;
      RECT 1.4600 1.0700 1.5500 1.3000 ;
      RECT 0.8600 1.3900 0.9500 1.6500 ;
      RECT 0.8600 0.8900 0.9500 1.3000 ;
      RECT 0.6000 0.8000 0.9500 0.8900 ;
      RECT 0.6000 0.4800 0.6900 0.8000 ;
  END
END AO22_X0P7M_A12TH

MACRO AO22_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 1.3950 0.3200 1.4950 0.4400 ;
        RECT 0.0800 0.3200 0.1700 0.7200 ;
        RECT 1.0850 0.4400 1.4950 0.5400 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0500 0.1600 1.4350 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4300 1.0500 0.5500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.7700 1.1500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 1.3700 1.7700 1.4600 2.0800 ;
        RECT 0.3400 1.7200 0.4300 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0100 0.7650 1.3600 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9700 1.7500 1.4350 ;
        RECT 1.6300 1.4350 1.7500 1.8650 ;
        RECT 1.6300 0.5600 1.7500 0.9700 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5400 0.6900 1.6300 ;
      RECT 0.6000 1.6300 0.6900 1.8300 ;
      RECT 0.6000 1.8300 1.2100 1.9200 ;
      RECT 1.1200 1.5100 1.2100 1.8300 ;
      RECT 0.0800 1.6300 0.1700 1.9600 ;
      RECT 0.8600 1.3000 1.5450 1.3900 ;
      RECT 1.4550 1.0300 1.5450 1.3000 ;
      RECT 0.8600 1.3900 0.9500 1.7100 ;
      RECT 0.8600 0.7150 0.9500 1.3000 ;
      RECT 0.5600 0.6250 0.9500 0.7150 ;
      RECT 0.5600 0.4250 0.7300 0.6250 ;
  END
END AO22_X1M_A12TH

MACRO AO22_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7050 ;
        RECT 1.1100 0.3200 1.2200 0.5200 ;
        RECT 2.1700 0.3200 2.5800 0.4500 ;
        RECT 3.0200 0.3200 3.1100 0.7200 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 1.2500 1.1150 1.3500 ;
        RECT 1.0150 0.8550 1.1150 1.2500 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0500 0.8850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2650 0.8500 2.2350 0.9500 ;
        RECT 1.2650 0.9500 1.3650 1.1600 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 0.3400 1.6750 0.4300 2.0800 ;
        RECT 0.8600 1.6750 0.9500 2.0800 ;
        RECT 2.5000 1.5950 2.5900 2.0800 ;
        RECT 3.0200 1.5950 3.1100 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5100 1.0500 1.9300 1.1600 ;
    END
    ANTENNAGATEAREA 0.1176 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9400 3.1500 1.2500 ;
        RECT 2.7550 1.2500 3.1500 1.3500 ;
        RECT 2.7550 0.8400 3.1500 0.9400 ;
        RECT 2.7550 1.3500 2.8550 1.8100 ;
        RECT 2.7550 0.4300 2.8550 0.8400 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 1.4800 1.2100 1.5700 ;
      RECT 1.1200 1.5700 1.2100 1.8300 ;
      RECT 1.1200 1.8300 2.2500 1.9200 ;
      RECT 1.6400 1.5100 1.7300 1.8300 ;
      RECT 2.1600 1.5100 2.2500 1.8300 ;
      RECT 0.0800 1.5700 0.1700 1.9100 ;
      RECT 0.6000 1.5700 0.6900 1.9100 ;
      RECT 2.4550 1.0550 2.9300 1.1450 ;
      RECT 1.3800 1.3000 2.5450 1.3900 ;
      RECT 2.4550 1.1450 2.5450 1.3000 ;
      RECT 2.4550 0.7000 2.5450 1.0550 ;
      RECT 0.6000 0.6100 2.5450 0.7000 ;
      RECT 1.9000 1.3900 1.9900 1.6500 ;
      RECT 1.6400 0.4850 1.7300 0.6100 ;
      RECT 1.3800 1.3900 1.4700 1.6500 ;
      RECT 0.6000 0.4850 0.6900 0.6100 ;
  END
END AO22_X1P4M_A12TH

MACRO AO22_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6700 ;
        RECT 1.0800 0.3200 1.2500 0.5450 ;
        RECT 2.1650 0.3200 2.5950 0.3900 ;
        RECT 3.0200 0.3200 3.1100 0.6700 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 0.8500 1.1150 0.9500 ;
        RECT 1.0150 0.9500 1.1150 1.2500 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0500 0.8850 1.1500 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2700 0.8500 2.2350 0.9500 ;
        RECT 1.2700 0.9500 1.3700 1.2200 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.2450 2.7200 ;
        RECT 2.5000 1.7700 2.5900 2.0800 ;
        RECT 3.0200 1.7700 3.1100 2.0800 ;
        RECT 0.3400 1.7200 0.4300 2.0800 ;
        RECT 0.8600 1.7200 0.9500 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5050 1.0500 1.9250 1.1500 ;
    END
    ANTENNAGATEAREA 0.1512 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9350 3.1500 1.3000 ;
        RECT 2.7550 1.3000 3.1500 1.4000 ;
        RECT 2.7550 0.8350 3.1500 0.9350 ;
        RECT 2.7550 1.4000 2.8550 1.7300 ;
        RECT 2.7550 0.5050 2.8550 0.8350 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5000 1.2100 1.5900 ;
      RECT 1.1200 1.5900 1.2100 1.8300 ;
      RECT 1.1200 1.8300 2.2500 1.9200 ;
      RECT 1.6400 1.5300 1.7300 1.8300 ;
      RECT 2.1600 1.5300 2.2500 1.8300 ;
      RECT 0.0800 1.5900 0.1700 1.9300 ;
      RECT 0.6000 1.5900 0.6900 1.9300 ;
      RECT 2.4550 1.0900 2.9300 1.1800 ;
      RECT 1.3800 1.3200 2.5450 1.4100 ;
      RECT 1.9000 1.4100 1.9900 1.7100 ;
      RECT 2.4550 1.1800 2.5450 1.3200 ;
      RECT 2.4550 0.7300 2.5450 1.0900 ;
      RECT 0.5600 0.6400 2.5450 0.7300 ;
      RECT 1.6000 0.4300 1.7700 0.6400 ;
      RECT 1.3800 1.4100 1.4700 1.7100 ;
      RECT 0.5600 0.4300 0.7300 0.6400 ;
  END
END AO22_X2M_A12TH

MACRO AO22_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6500 ;
        RECT 1.1200 0.3200 1.2100 0.4500 ;
        RECT 2.1600 0.3200 2.2500 0.4500 ;
        RECT 3.1650 0.3200 3.5750 0.3650 ;
        RECT 3.9700 0.3200 4.0600 0.6700 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 0.8500 1.3450 0.9500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4150 1.0500 1.5750 1.1500 ;
        RECT 1.4750 0.9350 1.5750 1.0500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9750 1.0500 3.2750 1.1500 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 3.4500 1.7700 3.5400 2.0800 ;
        RECT 3.9700 1.7700 4.0600 2.0800 ;
        RECT 0.3400 1.7150 0.4300 2.0800 ;
        RECT 0.8600 1.7150 0.9500 2.0800 ;
        RECT 1.3800 1.7150 1.4700 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7400 0.8500 2.9050 0.9500 ;
        RECT 1.7400 0.9500 1.8400 1.1450 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.9500 4.3500 1.3000 ;
        RECT 3.7050 1.3000 4.3500 1.4000 ;
        RECT 3.7050 0.8500 4.3500 0.9500 ;
        RECT 3.7050 1.4000 3.8050 1.7300 ;
        RECT 4.2300 1.4000 4.3500 1.7300 ;
        RECT 3.7050 0.5200 3.8050 0.8500 ;
        RECT 4.2300 0.5200 4.3500 0.8500 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5000 1.7300 1.5900 ;
      RECT 1.6400 1.5900 1.7300 1.8300 ;
      RECT 1.6400 1.8300 3.2900 1.9200 ;
      RECT 2.1600 1.5300 2.2500 1.8300 ;
      RECT 2.6800 1.5300 2.7700 1.8300 ;
      RECT 3.2000 1.5300 3.2900 1.8300 ;
      RECT 0.0800 1.5900 0.1700 1.9300 ;
      RECT 0.6000 1.5900 0.6900 1.9300 ;
      RECT 1.1200 1.5900 1.2100 1.9300 ;
      RECT 3.4800 1.0900 4.1050 1.1800 ;
      RECT 1.9000 1.4100 1.9900 1.7100 ;
      RECT 1.6000 0.4100 1.7700 0.6100 ;
      RECT 1.9000 1.3200 3.5700 1.4100 ;
      RECT 2.4200 1.4100 2.5100 1.7100 ;
      RECT 2.9400 1.4100 3.0300 1.7100 ;
      RECT 3.4800 1.1800 3.5700 1.3200 ;
      RECT 3.4800 0.7000 3.5700 1.0900 ;
      RECT 0.5600 0.6100 3.5700 0.7000 ;
      RECT 2.6400 0.4100 2.8100 0.6100 ;
      RECT 0.5600 0.4100 0.7300 0.6100 ;
  END
END AO22_X3M_A12TH

MACRO AO22_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6550 ;
        RECT 1.1200 0.3200 1.2100 0.4550 ;
        RECT 2.1600 0.3200 2.2500 0.4550 ;
        RECT 3.1900 0.3200 3.3000 0.4550 ;
        RECT 4.2550 0.3200 4.6550 0.3950 ;
        RECT 5.1050 0.3200 5.1950 0.6750 ;
        RECT 5.6250 0.3200 5.7150 0.6750 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.8500 2.1500 0.9500 ;
        RECT 0.2500 0.9500 0.3500 1.2500 ;
        RECT 2.0500 0.9500 2.1500 1.2500 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9400 5.7500 1.3000 ;
        RECT 4.8400 1.3000 5.7500 1.4000 ;
        RECT 4.8400 0.8400 5.7500 0.9400 ;
        RECT 4.8400 1.4000 4.9400 1.7300 ;
        RECT 5.3650 1.4000 5.4550 1.7300 ;
        RECT 4.8400 0.5100 4.9400 0.8400 ;
        RECT 5.3650 0.5050 5.4550 0.8400 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 4.5850 1.7700 4.6750 2.0800 ;
        RECT 5.1050 1.7700 5.1950 2.0800 ;
        RECT 5.6250 1.7700 5.7150 2.0800 ;
        RECT 0.3400 1.7200 0.4300 2.0800 ;
        RECT 0.8600 1.7200 0.9500 2.0800 ;
        RECT 1.3800 1.7200 1.4700 2.0800 ;
        RECT 1.9000 1.7200 1.9900 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5450 1.0500 3.9750 1.1500 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3050 0.8500 4.2300 0.9500 ;
        RECT 2.3050 0.9500 2.4050 1.2200 ;
        RECT 4.1300 0.9500 4.2300 1.2200 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.0500 1.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.3024 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5100 2.2500 1.6000 ;
      RECT 2.1600 1.6000 2.2500 1.8300 ;
      RECT 2.1600 1.8300 4.3300 1.9200 ;
      RECT 2.6800 1.5300 2.7700 1.8300 ;
      RECT 3.2000 1.5300 3.2900 1.8300 ;
      RECT 3.7200 1.5300 3.8100 1.8300 ;
      RECT 4.2400 1.5300 4.3300 1.8300 ;
      RECT 0.0800 1.6000 0.1700 1.9400 ;
      RECT 0.6000 1.6000 0.6900 1.9400 ;
      RECT 1.1200 1.6000 1.2100 1.9400 ;
      RECT 1.6400 1.6000 1.7300 1.9400 ;
      RECT 4.4800 1.0900 5.3600 1.1800 ;
      RECT 0.5600 0.4200 0.7300 0.6200 ;
      RECT 1.6000 0.4200 1.7700 0.6200 ;
      RECT 2.9400 1.4100 3.0300 1.7100 ;
      RECT 2.6400 0.4200 2.8100 0.6200 ;
      RECT 2.4200 1.4100 2.5100 1.7100 ;
      RECT 2.4200 1.3200 4.5700 1.4100 ;
      RECT 4.4800 1.1800 4.5700 1.3200 ;
      RECT 4.4800 0.7100 4.5700 1.0900 ;
      RECT 0.5600 0.6200 4.5700 0.7100 ;
      RECT 3.4600 1.4100 3.5500 1.7100 ;
      RECT 3.9800 1.4100 4.0700 1.7100 ;
      RECT 3.6800 0.4200 3.8500 0.6200 ;
  END
END AO22_X4M_A12TH

MACRO AO22_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.4450 0.3200 ;
        RECT 0.1000 0.3200 0.1900 0.6100 ;
        RECT 1.1000 0.3200 1.2700 0.5050 ;
        RECT 2.1400 0.3200 2.3100 0.5050 ;
        RECT 3.1800 0.3200 3.3500 0.5050 ;
        RECT 4.2200 0.3200 4.3900 0.5050 ;
        RECT 5.3150 0.3200 5.7250 0.3500 ;
        RECT 6.1700 0.3200 6.2600 0.6100 ;
        RECT 6.6900 0.3200 6.7800 0.6100 ;
        RECT 7.2100 0.3200 7.3000 0.6100 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9500 0.3500 1.1900 ;
        RECT 0.2500 0.8500 2.1350 0.9500 ;
        RECT 2.0350 0.9500 2.1350 1.0500 ;
        RECT 0.9850 0.9500 1.3950 1.0200 ;
        RECT 2.0350 1.0500 2.4200 1.1500 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0500 0.9150 7.1500 1.3000 ;
        RECT 5.9050 1.3000 7.1500 1.4000 ;
        RECT 5.9050 0.8150 7.1500 0.9150 ;
        RECT 5.9050 1.4000 6.0050 1.7300 ;
        RECT 6.4300 1.4000 6.5200 1.7300 ;
        RECT 6.9500 1.4000 7.0400 1.7300 ;
        RECT 5.9050 0.5050 6.0050 0.8150 ;
        RECT 6.4300 0.5050 6.5200 0.8150 ;
        RECT 6.9500 0.5050 7.0400 0.8150 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.4450 2.7200 ;
        RECT 0.3600 1.7850 0.4500 2.0800 ;
        RECT 0.8800 1.7850 0.9700 2.0800 ;
        RECT 1.4000 1.7850 1.4900 2.0800 ;
        RECT 1.9200 1.7850 2.0100 2.0800 ;
        RECT 2.4400 1.7850 2.5300 2.0800 ;
        RECT 5.6500 1.7700 5.7400 2.0800 ;
        RECT 6.1700 1.7700 6.2600 2.0800 ;
        RECT 6.6900 1.7700 6.7800 2.0800 ;
        RECT 7.2100 1.7700 7.3000 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.8500 5.0550 0.9500 ;
        RECT 2.8500 0.9500 2.9500 1.1450 ;
        RECT 3.6050 0.9500 4.0050 1.0150 ;
        RECT 4.6450 0.9500 5.0550 1.0100 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0800 1.0500 3.4700 1.1300 ;
        RECT 3.0800 1.1300 5.3500 1.2300 ;
        RECT 4.1200 1.0500 4.5100 1.1300 ;
        RECT 5.2500 0.9350 5.3500 1.1300 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END B1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 2.6450 1.3500 ;
        RECT 0.7700 1.1500 0.8700 1.2500 ;
        RECT 1.5250 1.1500 1.6250 1.2500 ;
        RECT 2.5450 0.9350 2.6450 1.2500 ;
        RECT 0.4750 1.0500 0.8700 1.1500 ;
        RECT 1.5250 1.0500 1.9150 1.1500 ;
    END
    ANTENNAGATEAREA 0.4485 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.1000 1.5000 2.7900 1.5900 ;
      RECT 2.7000 1.5900 2.7900 1.8300 ;
      RECT 2.7000 1.8300 5.3900 1.9200 ;
      RECT 3.2200 1.5300 3.3100 1.8300 ;
      RECT 3.7400 1.5300 3.8300 1.8300 ;
      RECT 4.2600 1.5300 4.3500 1.8300 ;
      RECT 4.7800 1.5300 4.8700 1.8300 ;
      RECT 5.3000 1.5300 5.3900 1.8300 ;
      RECT 0.1000 1.5900 0.1900 1.9500 ;
      RECT 0.6200 1.5900 0.7100 1.9100 ;
      RECT 1.1400 1.5900 1.2300 1.9300 ;
      RECT 1.6600 1.5900 1.7500 1.9300 ;
      RECT 2.1800 1.5900 2.2700 1.9300 ;
      RECT 5.6550 1.0900 6.8050 1.1800 ;
      RECT 0.5800 0.4300 0.7500 0.6300 ;
      RECT 1.6200 0.4300 1.7900 0.6300 ;
      RECT 2.6600 0.4300 2.8300 0.6300 ;
      RECT 2.9600 1.4100 3.0500 1.7100 ;
      RECT 3.4800 1.4100 3.5700 1.7100 ;
      RECT 4.0000 1.4100 4.0900 1.7100 ;
      RECT 3.7000 0.4300 3.8700 0.6300 ;
      RECT 2.9600 1.3200 5.7450 1.4100 ;
      RECT 5.6550 1.1800 5.7450 1.3200 ;
      RECT 5.6550 0.7200 5.7450 1.0900 ;
      RECT 0.5800 0.6300 5.7450 0.7200 ;
      RECT 5.0400 1.4100 5.1300 1.7100 ;
      RECT 4.7400 0.4300 4.9100 0.6300 ;
      RECT 4.5200 1.4100 4.6100 1.7100 ;
  END
END AO22_X6M_A12TH

MACRO AOI211_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6150 0.3200 0.7850 0.5100 ;
        RECT 1.1400 0.3200 1.3100 0.5100 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9900 0.3500 1.4100 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3800 1.7600 0.4800 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9900 0.5600 1.4100 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7750 0.8100 0.9500 1.1000 ;
    END
    ANTENNAGATEAREA 0.0348 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.9900 1.1500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0348 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.5500 ;
        RECT 1.1750 1.5500 1.3500 1.6500 ;
        RECT 0.1200 0.6000 1.3500 0.7000 ;
        RECT 1.1750 1.6500 1.2750 1.9600 ;
        RECT 0.8800 0.4250 1.0500 0.6000 ;
        RECT 0.1200 0.4100 0.2200 0.6000 ;
    END
    ANTENNADIFFAREA 0.15825 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5400 0.7500 1.6400 ;
      RECT 0.6500 1.6400 0.7500 1.9700 ;
      RECT 0.1200 1.6400 0.2200 1.9700 ;
  END
END AOI211_X0P5M_A12TH

MACRO AOI211_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6150 0.3200 0.7850 0.5100 ;
        RECT 1.1400 0.3200 1.3100 0.5100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3800 1.7000 0.4800 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.5000 ;
        RECT 1.1750 1.5000 1.3500 1.6000 ;
        RECT 0.1200 0.6000 1.3500 0.7000 ;
        RECT 1.1750 1.6000 1.2750 1.9300 ;
        RECT 0.1200 0.4850 0.2200 0.6000 ;
        RECT 0.9150 0.4150 1.0150 0.6000 ;
    END
    ANTENNADIFFAREA 0.2236 ;
  END Y

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.9350 1.1500 1.3250 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.9350 0.8400 1.3900 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END B0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9350 0.5600 1.3750 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9350 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0552 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5000 0.7500 1.6000 ;
      RECT 0.6500 1.6000 0.7500 1.9300 ;
      RECT 0.1200 1.6000 0.2200 1.9300 ;
  END
END AOI211_X0P7M_A12TH

MACRO AOI211_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6400 0.3200 0.7400 0.5100 ;
        RECT 1.1750 0.3200 1.2750 0.5100 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3800 1.7700 0.4800 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0400 0.1600 1.4250 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.7900 0.5600 1.1600 ;
    END
    ANTENNAGATEAREA 0.078 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 0.8050 0.9500 1.0300 ;
        RECT 0.7100 1.0300 0.9500 1.1200 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 0.8650 1.1500 1.3200 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END C0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7000 1.3500 1.5150 ;
        RECT 1.1750 1.5150 1.3500 1.6150 ;
        RECT 0.0850 0.6000 1.3500 0.7000 ;
        RECT 1.1750 1.6150 1.2750 1.9450 ;
        RECT 0.0850 0.4100 0.2550 0.6000 ;
        RECT 0.9150 0.4100 1.0150 0.6000 ;
    END
    ANTENNADIFFAREA 0.3165 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.1200 1.5150 0.7500 1.6150 ;
      RECT 0.6500 1.6150 0.7500 1.9450 ;
      RECT 0.1200 1.6150 0.2200 1.9450 ;
  END
END AOI211_X1M_A12TH

MACRO AOI211_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.3000 1.6500 0.4700 2.0800 ;
        RECT 0.8200 1.6500 0.9900 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.5600 ;
        RECT 1.1150 0.3200 1.2150 0.5600 ;
        RECT 1.6450 0.3200 1.7450 0.5600 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1400 1.0500 1.1200 1.1500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.8500 0.9200 0.9500 ;
    END
    ANTENNAGATEAREA 0.1104 ;
  END A0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4800 1.0500 1.9000 1.1750 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1950 0.8500 1.9250 0.9500 ;
    END
    ANTENNAGATEAREA 0.0984 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.7500 2.1500 1.3000 ;
        RECT 1.5750 1.3000 2.1500 1.4000 ;
        RECT 0.5950 0.6500 2.1500 0.7500 ;
        RECT 1.5750 1.4000 1.6750 1.6900 ;
        RECT 1.3850 0.5150 1.4850 0.6500 ;
        RECT 0.5950 0.4400 0.6950 0.6500 ;
    END
    ANTENNADIFFAREA 0.254 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.1200 1.7900 2.1250 1.8900 ;
      RECT 2.0250 1.5200 2.1250 1.7900 ;
      RECT 0.0750 1.4600 1.2200 1.5600 ;
      RECT 1.1200 1.5600 1.2200 1.7900 ;
      RECT 0.0750 1.5600 0.1750 1.9100 ;
      RECT 0.5950 1.5600 0.6950 1.9100 ;
  END
END AOI211_X1P4M_A12TH

MACRO AOI211_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0850 0.3200 0.2550 0.6700 ;
        RECT 1.1700 0.3200 1.2700 0.5600 ;
        RECT 1.6700 0.3200 1.8400 0.5600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3800 1.7700 0.4800 2.0800 ;
        RECT 0.9000 1.7700 1.0000 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.7500 2.3500 1.2800 ;
        RECT 1.6800 1.2800 2.3500 1.3800 ;
        RECT 0.6050 0.6500 2.3500 0.7500 ;
        RECT 1.6800 1.3800 1.7800 1.7000 ;
        RECT 0.6050 0.4350 0.7750 0.6500 ;
        RECT 1.4000 0.4350 1.5700 0.6500 ;
    END
    ANTENNADIFFAREA 0.365 ;
  END Y

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2600 0.8500 2.1250 0.9500 ;
        RECT 1.2600 0.9500 1.3600 1.1300 ;
        RECT 2.0250 0.9500 2.1250 1.1400 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END B0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4800 1.0500 1.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.1392 ;
  END C0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 0.8850 1.1500 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2500 1.1050 1.3500 ;
        RECT 0.2500 1.1550 0.3500 1.2500 ;
        RECT 1.0050 1.0400 1.1050 1.2500 ;
        RECT 0.0850 1.0550 0.3500 1.1550 ;
    END
    ANTENNAGATEAREA 0.156 ;
  END A1
  OBS
    LAYER M1 ;
      RECT 1.1700 1.8100 2.2800 1.9100 ;
      RECT 2.1800 1.5200 2.2800 1.8100 ;
      RECT 0.1200 1.4800 1.2700 1.5800 ;
      RECT 1.1700 1.5800 1.2700 1.8100 ;
      RECT 0.1200 1.5800 0.2200 1.9100 ;
      RECT 0.6400 1.5800 0.7400 1.9100 ;
  END
END AOI211_X2M_A12TH

MACRO AOI211_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.8100 ;
        RECT 1.1300 0.3200 1.2300 0.5600 ;
        RECT 1.9100 0.3200 2.0100 0.5600 ;
        RECT 2.4300 0.3200 2.5300 0.5600 ;
        RECT 2.9500 0.3200 3.0500 0.5600 ;
    END
  END VSS

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6400 1.0500 3.1100 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END C0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.3500 1.7700 0.4500 2.0800 ;
        RECT 0.8700 1.7700 0.9700 2.0800 ;
        RECT 1.3900 1.7700 1.4900 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8550 1.0450 2.3200 1.1500 ;
    END
    ANTENNAGATEAREA 0.2088 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.7500 3.3500 1.3000 ;
        RECT 2.6900 1.3000 3.3500 1.4000 ;
        RECT 0.5750 0.6500 3.3500 0.7500 ;
        RECT 2.6900 1.4000 2.7900 1.7000 ;
        RECT 3.2100 1.4000 3.3500 1.7200 ;
        RECT 1.6250 0.4400 1.7250 0.6500 ;
        RECT 2.1700 0.4400 2.2700 0.6500 ;
        RECT 2.6900 0.4400 2.7900 0.6500 ;
        RECT 3.2100 0.4400 3.3100 0.6500 ;
        RECT 0.5750 0.4200 0.7450 0.6500 ;
    END
    ANTENNADIFFAREA 0.6416 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.2900 1.1500 1.3900 ;
        RECT 1.0500 1.1500 1.1500 1.2900 ;
        RECT 0.2500 1.1450 0.3500 1.2900 ;
        RECT 1.0500 1.0500 1.3300 1.1500 ;
        RECT 0.1200 1.0550 0.3500 1.1450 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4750 1.0500 0.8500 1.1500 ;
        RECT 0.7500 0.9500 0.8500 1.0500 ;
        RECT 0.7500 0.8500 1.6000 0.9500 ;
        RECT 1.5000 0.9500 1.6000 1.1200 ;
    END
    ANTENNAGATEAREA 0.234 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0900 1.5000 2.2700 1.6000 ;
      RECT 1.6500 1.6000 1.7500 1.9300 ;
      RECT 2.1700 1.6000 2.2700 1.7100 ;
      RECT 0.0900 1.6000 0.1900 1.9300 ;
      RECT 0.6100 1.6000 0.7100 1.9300 ;
      RECT 1.1300 1.6000 1.2300 1.9300 ;
      RECT 1.9100 1.8200 3.0500 1.9200 ;
      RECT 2.9500 1.5100 3.0500 1.8200 ;
      RECT 1.9100 1.7100 2.0100 1.8200 ;
      RECT 2.4300 1.4900 2.5300 1.8200 ;
  END
END AOI211_X3M_A12TH

MACRO AOI211_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 1.1300 0.3200 1.2300 0.5100 ;
        RECT 2.1450 0.3200 2.2450 0.5100 ;
        RECT 2.6900 0.3200 2.7900 0.5100 ;
        RECT 3.2100 0.3200 3.3100 0.5100 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9750 1.0500 1.3900 1.1500 ;
        RECT 0.9750 1.1500 1.0750 1.2500 ;
        RECT 0.2450 1.2500 2.1150 1.3500 ;
        RECT 0.2450 1.1800 0.3450 1.2500 ;
        RECT 2.0150 1.0400 2.1150 1.2500 ;
        RECT 0.0950 1.0800 0.3450 1.1800 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4750 1.0500 0.8500 1.1500 ;
        RECT 0.7500 0.9500 0.8500 1.0500 ;
        RECT 0.7500 0.8500 1.6150 0.9500 ;
        RECT 1.5150 0.9500 1.6150 1.0500 ;
        RECT 1.5150 1.0500 1.8900 1.1500 ;
    END
    ANTENNAGATEAREA 0.312 ;
  END A0

  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5550 1.0500 2.9300 1.1500 ;
        RECT 2.8300 0.9500 2.9300 1.0500 ;
        RECT 2.8300 0.8500 3.7050 0.9500 ;
        RECT 3.5750 0.9500 3.7050 1.0500 ;
        RECT 3.5750 1.0500 3.9450 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END C0

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2900 1.2500 4.1550 1.3500 ;
        RECT 2.2900 1.1500 2.4100 1.2500 ;
        RECT 3.0400 1.1500 3.1400 1.2500 ;
        RECT 4.0550 0.9250 4.1550 1.2500 ;
        RECT 2.2400 1.0600 2.4100 1.1500 ;
        RECT 3.0400 1.0500 3.4500 1.1500 ;
    END
    ANTENNAGATEAREA 0.2784 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2500 0.7200 4.3500 1.4400 ;
        RECT 2.6550 1.4400 4.3500 1.5400 ;
        RECT 0.5750 0.6200 4.3500 0.7200 ;
        RECT 2.6550 1.5400 2.8250 1.7300 ;
        RECT 3.6750 1.5400 3.8450 1.7300 ;
        RECT 0.5750 0.4100 0.7450 0.6200 ;
        RECT 1.6150 0.4100 1.7850 0.6200 ;
        RECT 2.3950 0.4100 2.5650 0.6200 ;
        RECT 2.9150 0.4100 3.0850 0.6200 ;
    END
    ANTENNADIFFAREA 0.7746 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 0.3500 1.7900 0.4500 2.0800 ;
        RECT 0.8700 1.7900 0.9700 2.0800 ;
        RECT 1.3900 1.7900 1.4900 2.0800 ;
        RECT 1.9100 1.7900 2.0100 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1700 1.8200 4.3500 1.9200 ;
      RECT 4.1750 1.6300 4.3450 1.8200 ;
      RECT 2.1700 1.6000 2.2700 1.8200 ;
      RECT 0.0900 1.5000 2.2700 1.6000 ;
      RECT 0.0900 1.6000 0.1900 1.9100 ;
      RECT 0.6100 1.6000 0.7100 1.9100 ;
      RECT 1.1300 1.6000 1.2300 1.9100 ;
      RECT 1.6500 1.6000 1.7500 1.9100 ;
      RECT 3.1750 1.6300 3.3450 1.8200 ;
  END
END AOI211_X4M_A12TH

MACRO AOI21B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1800 0.5200 ;
        RECT 0.9450 0.3200 1.0350 0.6300 ;
        RECT 1.2300 0.3200 1.3200 0.9100 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2450 0.9000 0.3500 1.3000 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.6950 0.5500 1.1150 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0050 1.0350 1.3500 1.1600 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END B0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8400 1.6100 1.0100 1.9900 ;
        RECT 0.7500 1.5500 1.0100 1.6100 ;
        RECT 0.6400 1.5200 1.0100 1.5500 ;
        RECT 0.6400 1.4500 0.8400 1.5200 ;
        RECT 0.6400 0.4600 0.7300 1.4500 ;
    END
    ANTENNADIFFAREA 0.1408 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3100 1.8200 0.4800 2.0800 ;
        RECT 1.2300 1.3000 1.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.7000 0.7500 1.7300 ;
      RECT 0.5700 1.7300 0.7500 1.9900 ;
      RECT 0.0500 1.6400 0.6600 1.7000 ;
      RECT 0.0500 1.7300 0.2200 1.9900 ;
      RECT 0.9300 1.3600 1.1000 1.4100 ;
      RECT 0.8250 1.2700 1.1000 1.3600 ;
      RECT 0.8250 0.8350 1.0600 0.9250 ;
      RECT 0.9700 0.7200 1.0600 0.8350 ;
      RECT 0.8250 0.9250 0.9150 1.2700 ;
  END
END AOI21B_X0P5M_A12TH

MACRO AOI21B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6300 ;
        RECT 0.8800 0.3200 0.9900 0.4600 ;
        RECT 1.4100 0.3200 1.5100 0.6350 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9500 0.5500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.7750 0.1600 1.1700 ;
    END
    ANTENNAGATEAREA 0.0639 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 0.8150 1.5500 1.2150 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END B0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3500 1.7400 0.4500 2.0800 ;
        RECT 1.4100 1.4100 1.5100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.7500 0.9500 1.5250 ;
        RECT 0.8500 1.5250 1.0200 1.9350 ;
        RECT 0.5600 0.6500 0.9500 0.7500 ;
        RECT 0.5600 0.4300 0.6600 0.6500 ;
    END
    ANTENNADIFFAREA 0.203925 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5300 0.7050 1.6200 ;
      RECT 0.6150 1.6200 0.7050 1.9600 ;
      RECT 0.0950 1.6200 0.1850 1.9600 ;
      RECT 1.1550 1.4200 1.2450 1.6300 ;
      RECT 1.0650 1.3300 1.2450 1.4200 ;
      RECT 1.0650 0.7200 1.1550 1.3300 ;
      RECT 1.0650 0.6300 1.2450 0.7200 ;
      RECT 1.1550 0.4400 1.2450 0.6300 ;
  END
END AOI21B_X0P7M_A12TH

MACRO AOI21B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.0850 0.3200 0.1750 0.8900 ;
        RECT 0.5900 0.3200 0.6900 0.9250 ;
        RECT 1.4100 0.3200 1.5100 0.7350 ;
    END
  END VSS

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0100 0.1650 1.4300 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END B0N

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9700 1.1500 1.3950 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4400 0.9350 1.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.09 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.4900 0.9500 1.2900 ;
        RECT 0.5900 1.2900 0.9500 1.3900 ;
        RECT 0.5900 1.3900 0.6900 1.7200 ;
    END
    ANTENNADIFFAREA 0.260325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 1.1500 1.7700 1.2500 2.0800 ;
        RECT 0.0800 1.5500 0.1800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3400 1.0450 0.7300 1.1550 ;
      RECT 0.3400 1.1550 0.4400 1.7450 ;
      RECT 0.3400 0.6950 0.4400 1.0450 ;
      RECT 0.8450 1.5200 1.5150 1.6200 ;
      RECT 1.4050 1.6200 1.5150 1.9500 ;
      RECT 0.8450 1.6200 0.9550 1.9500 ;
  END
END AOI21B_X1M_A12TH

MACRO AOI21B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.8250 ;
        RECT 1.1300 0.3200 1.2300 0.6150 ;
        RECT 1.7100 0.3200 1.8100 0.6150 ;
        RECT 2.2200 0.3200 2.3200 0.7950 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.4600 1.5500 0.8500 ;
        RECT 0.6100 0.8500 1.5500 0.9500 ;
        RECT 1.2500 0.9500 1.3500 1.2800 ;
        RECT 0.6100 0.4350 0.7100 0.8500 ;
        RECT 1.2500 1.2800 1.4900 1.3800 ;
        RECT 1.3900 1.3800 1.4900 1.7050 ;
    END
    ANTENNADIFFAREA 0.266 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.3500 1.7300 0.4500 2.0800 ;
        RECT 0.8700 1.7300 0.9700 2.0800 ;
        RECT 2.2250 1.6650 2.3250 2.0800 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2500 1.1500 1.3500 ;
        RECT 1.0500 1.0850 1.1500 1.2500 ;
        RECT 0.0500 0.9850 0.1600 1.2500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0500 0.8650 1.1500 ;
    END
    ANTENNAGATEAREA 0.1278 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9000 1.0500 2.3300 1.1500 ;
    END
    ANTENNAGATEAREA 0.0333 ;
  END B0N
  OBS
    LAYER M1 ;
      RECT 1.1300 1.8200 1.7500 1.9200 ;
      RECT 1.6500 1.5100 1.7500 1.8200 ;
      RECT 0.0900 1.5050 1.2300 1.6050 ;
      RECT 1.1300 1.6050 1.2300 1.8200 ;
      RECT 0.0900 1.6050 0.1900 1.9550 ;
      RECT 0.6100 1.6050 0.7100 1.9550 ;
      RECT 1.9600 1.3900 2.0600 1.7800 ;
      RECT 1.6500 1.2900 2.0600 1.3900 ;
      RECT 1.6500 0.8500 2.0600 0.9500 ;
      RECT 1.9600 0.6250 2.0600 0.8500 ;
      RECT 1.6500 1.1550 1.7500 1.2900 ;
      RECT 1.5050 1.0550 1.7500 1.1550 ;
      RECT 1.6500 0.9500 1.7500 1.0550 ;
  END
END AOI21B_X1P4M_A12TH

MACRO AND4_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 1.0400 0.3200 1.1400 0.6700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9200 1.5500 1.4150 ;
        RECT 1.4050 1.4150 1.5500 1.5150 ;
        RECT 1.4050 0.8200 1.5500 0.9200 ;
        RECT 1.4050 1.5150 1.5050 1.8250 ;
        RECT 1.4050 0.5100 1.5050 0.8200 ;
    END
    ANTENNADIFFAREA 0.202125 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9700 0.5600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.4500 0.9050 1.5500 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.0500 1.1150 1.1500 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9700 0.1600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0579 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.0900 1.8500 0.1900 2.0800 ;
        RECT 0.6100 1.8500 0.7100 2.0800 ;
        RECT 1.1450 1.8500 1.2450 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 1.6700 1.3000 1.7600 ;
      RECT 1.2100 1.2550 1.3000 1.6700 ;
      RECT 1.2100 1.0850 1.3450 1.2550 ;
      RECT 1.2100 0.8800 1.3000 1.0850 ;
      RECT 0.1300 0.7900 1.3000 0.8800 ;
      RECT 0.3550 1.7600 0.4450 1.9650 ;
      RECT 0.1300 0.4450 0.2200 0.7900 ;
      RECT 0.8750 1.7600 0.9650 1.9650 ;
  END
END AND4_X0P7M_A12TH

MACRO AND4_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 1.3000 0.3200 1.4700 0.5300 ;
        RECT 1.7200 0.3200 1.8900 0.5300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 1.7550 1.7700 1.8550 2.0800 ;
        RECT 0.8200 1.7550 0.9900 2.0800 ;
        RECT 1.3400 1.7550 1.5100 2.0800 ;
        RECT 0.3350 1.6500 0.4350 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9200 2.1500 1.3100 ;
        RECT 2.0150 1.3100 2.1500 1.4100 ;
        RECT 2.0150 0.8200 2.1500 0.9200 ;
        RECT 2.0150 1.4100 2.1150 1.7400 ;
        RECT 2.0150 0.4900 2.1150 0.8200 ;
    END
    ANTENNADIFFAREA 0.27625 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5600 1.2800 ;
        RECT 0.2800 1.2800 0.5600 1.4300 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9650 1.2950 1.1500 1.4650 ;
        RECT 1.0500 1.0400 1.1500 1.2950 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.0800 0.7500 1.3650 ;
        RECT 0.6500 1.3650 0.8650 1.4550 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2800 1.2500 1.5900 1.4350 ;
    END
    ANTENNAGATEAREA 0.0912 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.5950 1.5650 1.8750 1.6650 ;
      RECT 1.7750 0.7200 1.8750 1.5650 ;
      RECT 1.1100 0.6200 1.8750 0.7200 ;
      RECT 0.5950 1.6650 0.6950 1.9700 ;
      RECT 0.3750 0.5800 0.4750 0.8700 ;
      RECT 1.1150 1.6650 1.2150 1.9900 ;
      RECT 1.1100 0.5800 1.2100 0.6200 ;
      RECT 0.3750 0.4800 1.2100 0.5800 ;
  END
END AND4_X1M_A12TH

MACRO AND4_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6500 ;
        RECT 1.8950 0.3200 1.9850 0.7350 ;
        RECT 2.4300 0.3200 2.5200 0.7850 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1700 1.2500 2.5550 1.3500 ;
        RECT 2.1700 1.3500 2.2600 1.9450 ;
        RECT 2.4650 0.9800 2.5550 1.2500 ;
        RECT 2.1700 0.8900 2.5550 0.9800 ;
        RECT 2.1700 0.4550 2.2600 0.8900 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 1.4700 1.7400 1.5300 ;
        RECT 0.8100 1.5300 0.9900 1.5500 ;
        RECT 0.8100 1.4400 1.8300 1.4700 ;
        RECT 0.8100 1.5500 0.9000 1.5950 ;
        RECT 1.6500 1.3800 1.8300 1.4400 ;
        RECT 0.2200 1.5950 0.9000 1.6850 ;
        RECT 1.7400 1.2600 1.8300 1.3800 ;
        RECT 0.2200 1.4750 0.3100 1.5950 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 0.8500 1.3900 0.9500 ;
        RECT 1.3000 0.9500 1.3900 1.0050 ;
        RECT 0.4000 0.9500 0.4900 1.3550 ;
        RECT 1.3000 1.0050 1.5900 1.0950 ;
        RECT 1.5000 1.0950 1.5900 1.2150 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.2500 1.4000 1.3500 ;
        RECT 0.6100 1.3500 0.7200 1.4850 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.0500 1.1900 1.1500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 0.8150 1.8400 0.9850 2.0800 ;
        RECT 1.3750 1.8000 1.4650 2.0800 ;
        RECT 1.9100 1.8000 2.0000 2.0800 ;
        RECT 2.4300 1.7300 2.5200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.9200 1.0700 2.3550 1.1600 ;
      RECT 1.1150 1.6200 2.0100 1.7100 ;
      RECT 1.9200 1.1600 2.0100 1.6200 ;
      RECT 1.9200 0.9150 2.0100 1.0700 ;
      RECT 1.4800 0.8250 2.0100 0.9150 ;
      RECT 1.1150 1.7100 1.2050 1.9900 ;
      RECT 0.9000 0.4700 1.0700 0.6700 ;
      RECT 1.4800 0.7600 1.5700 0.8250 ;
      RECT 0.9000 0.6700 1.5700 0.7600 ;
      RECT 1.6350 1.7100 1.7250 1.9900 ;
  END
END AND4_X1P4M_A12TH

MACRO AND4_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.6450 0.3200 ;
        RECT 0.9200 0.3200 1.0200 0.6300 ;
        RECT 2.8900 0.3200 2.9900 0.6350 ;
        RECT 3.4100 0.3200 3.5100 0.6350 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6900 1.2500 1.1550 1.3800 ;
    END
    ANTENNAGATEAREA 0.1572 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8100 1.2500 2.2300 1.3500 ;
    END
    ANTENNAGATEAREA 0.1572 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5950 1.0500 2.5800 1.1500 ;
        RECT 1.5950 1.1500 1.6950 1.3850 ;
        RECT 2.4800 1.1500 2.5800 1.3900 ;
    END
    ANTENNAGATEAREA 0.1572 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.0500 1.3850 1.1500 ;
        RECT 0.4000 1.1500 0.5000 1.3950 ;
        RECT 1.2850 1.1500 1.3850 1.3850 ;
    END
    ANTENNAGATEAREA 0.1572 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.9050 3.5500 1.2900 ;
        RECT 3.1500 1.2900 3.5500 1.3900 ;
        RECT 3.1500 0.8050 3.5500 0.9050 ;
        RECT 3.1500 1.3900 3.2500 1.7400 ;
        RECT 3.1500 0.4700 3.2500 0.8050 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.6450 2.7200 ;
        RECT 2.8900 1.7700 2.9900 2.0800 ;
        RECT 3.4100 1.7700 3.5100 2.0800 ;
        RECT 0.8850 1.6900 1.0550 2.0800 ;
        RECT 1.4050 1.6900 1.5750 2.0800 ;
        RECT 1.9250 1.6900 2.0950 2.0800 ;
        RECT 2.4450 1.6900 2.6150 2.0800 ;
        RECT 0.4050 1.5850 0.4950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.8550 1.0550 3.2900 1.1450 ;
      RECT 0.6650 1.4850 2.9450 1.5750 ;
      RECT 2.8550 1.1450 2.9450 1.4850 ;
      RECT 2.8550 0.9600 2.9450 1.0550 ;
      RECT 1.9250 0.8700 2.9450 0.9600 ;
      RECT 0.6650 1.5750 0.7550 1.9700 ;
      RECT 1.1850 1.5750 1.2750 1.9700 ;
      RECT 2.2250 1.5750 2.3150 1.9700 ;
      RECT 1.9250 0.6700 2.0950 0.8700 ;
      RECT 1.7050 1.5750 1.7950 1.9700 ;
      RECT 0.4050 0.8700 1.5350 0.9600 ;
      RECT 1.4450 0.5700 1.5350 0.8700 ;
      RECT 1.4450 0.4800 2.5750 0.5700 ;
      RECT 2.4850 0.5700 2.5750 0.7800 ;
      RECT 2.4850 0.4100 2.5750 0.4800 ;
      RECT 0.4050 0.5050 0.4950 0.8700 ;
  END
END AND4_X2M_A12TH

MACRO AND4_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.4650 0.3200 0.5650 0.6300 ;
        RECT 0.9850 0.3200 1.0850 0.6300 ;
        RECT 4.0300 0.3200 4.1300 0.6350 ;
        RECT 4.5500 0.3200 4.6500 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 4.0300 1.7700 4.1300 2.0800 ;
        RECT 4.5500 1.7700 4.6500 2.0800 ;
        RECT 1.2450 1.6850 1.3450 2.0800 ;
        RECT 1.7650 1.6850 1.8650 2.0800 ;
        RECT 2.2850 1.6850 2.3850 2.0800 ;
        RECT 2.8050 1.6850 2.9050 2.0800 ;
        RECT 3.3250 1.6850 3.4250 2.0800 ;
        RECT 0.7250 1.6450 0.8250 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.9500 4.9500 1.2500 ;
        RECT 4.2900 1.2500 4.9500 1.3500 ;
        RECT 4.2900 0.8500 4.9500 0.9500 ;
        RECT 4.2900 1.3500 4.3900 1.7350 ;
        RECT 4.8100 1.3500 4.9100 1.7350 ;
        RECT 4.2900 0.4750 4.3900 0.8500 ;
        RECT 4.8100 0.4750 4.9100 0.8500 ;
    END
    ANTENNADIFFAREA 0.609375 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4450 1.2500 1.9550 1.3500 ;
    END
    ANTENNAGATEAREA 0.2208 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2400 1.2500 2.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.2208 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0400 1.2500 3.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.2208 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.2500 1.1600 1.3500 ;
    END
    ANTENNAGATEAREA 0.2208 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.7300 0.8700 1.3400 0.9600 ;
      RECT 1.2500 0.5700 1.3400 0.8700 ;
      RECT 1.2500 0.4800 1.8600 0.5700 ;
      RECT 1.7700 0.5700 1.8600 0.9150 ;
      RECT 0.7300 0.5300 0.8200 0.8700 ;
      RECT 1.5100 1.0050 2.1150 1.0950 ;
      RECT 2.0250 0.9550 2.1150 1.0050 ;
      RECT 1.5100 0.6600 1.6000 1.0050 ;
      RECT 2.0250 0.5700 2.1200 0.9550 ;
      RECT 2.0250 0.4800 2.6400 0.5700 ;
      RECT 2.5500 0.5700 2.6400 0.9150 ;
      RECT 2.2900 1.0050 2.9000 1.0950 ;
      RECT 2.2900 0.6600 2.3800 1.0050 ;
      RECT 2.8100 0.5700 2.9000 1.0050 ;
      RECT 2.8100 0.4800 3.4200 0.5700 ;
      RECT 3.3300 0.5700 3.4200 0.8900 ;
      RECT 4.0550 1.1000 4.7050 1.1550 ;
      RECT 3.0700 1.0550 4.7050 1.1000 ;
      RECT 0.9900 1.5900 1.0800 1.9250 ;
      RECT 1.5100 1.5900 1.6000 1.9250 ;
      RECT 2.5500 1.5900 2.6400 1.9250 ;
      RECT 3.0700 1.5900 3.1600 1.9250 ;
      RECT 3.0700 0.6600 3.1600 1.0100 ;
      RECT 3.5850 0.6100 3.6850 1.0100 ;
      RECT 0.9900 1.5000 4.1450 1.5900 ;
      RECT 4.0550 1.1550 4.1450 1.5000 ;
      RECT 3.0700 1.0100 4.1450 1.0550 ;
  END
END AND4_X3M_A12TH

MACRO AND4_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.3650 0.3200 0.4550 0.6250 ;
        RECT 0.8850 0.3200 0.9750 0.6250 ;
        RECT 4.8250 0.3200 4.9250 0.6300 ;
        RECT 5.3450 0.3200 5.4450 0.6300 ;
        RECT 5.8650 0.3200 5.9650 0.6300 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3150 1.2500 1.0250 1.3500 ;
    END
    ANTENNAGATEAREA 0.306 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7250 1.2500 4.4350 1.3500 ;
    END
    ANTENNAGATEAREA 0.306 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7250 1.2500 3.4350 1.3500 ;
        RECT 2.7250 1.2450 2.8300 1.2500 ;
    END
    ANTENNAGATEAREA 0.306 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3350 1.2500 2.0450 1.3500 ;
    END
    ANTENNAGATEAREA 0.306 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9000 5.7500 1.3000 ;
        RECT 5.0850 1.3000 5.7500 1.4000 ;
        RECT 5.0850 0.8000 5.7500 0.9000 ;
        RECT 5.0850 1.4000 5.1850 1.7300 ;
        RECT 5.6050 1.4000 5.7050 1.7300 ;
        RECT 5.0850 0.4700 5.1850 0.8000 ;
        RECT 5.6050 0.4700 5.7050 0.8000 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 4.8250 1.7650 4.9250 2.0800 ;
        RECT 5.3450 1.7650 5.4450 2.0800 ;
        RECT 5.8650 1.7650 5.9650 2.0800 ;
        RECT 0.6250 1.7200 0.7150 2.0800 ;
        RECT 1.1450 1.7200 1.2350 2.0800 ;
        RECT 1.6650 1.7200 1.7550 2.0800 ;
        RECT 2.1850 1.7200 2.2750 2.0800 ;
        RECT 2.4650 1.7200 2.5550 2.0800 ;
        RECT 2.9850 1.7200 3.0750 2.0800 ;
        RECT 3.5050 1.7200 3.5950 2.0800 ;
        RECT 4.0250 1.7200 4.1150 2.0800 ;
        RECT 4.5450 1.7200 4.6350 2.0800 ;
        RECT 0.1050 1.5200 0.1950 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.1050 0.8650 1.2350 0.9550 ;
      RECT 1.1450 0.5700 1.2350 0.8650 ;
      RECT 1.1450 0.4800 2.2750 0.5700 ;
      RECT 1.6650 0.5700 1.7550 0.8850 ;
      RECT 2.1850 0.5700 2.2750 0.8850 ;
      RECT 0.1050 0.5250 0.1950 0.8650 ;
      RECT 0.6250 0.5250 0.7150 0.8650 ;
      RECT 1.4050 1.0000 3.3350 1.0900 ;
      RECT 1.4050 0.6800 1.4950 1.0000 ;
      RECT 1.9250 0.6800 2.0150 1.0000 ;
      RECT 2.7250 0.6800 2.8150 1.0000 ;
      RECT 3.2450 0.6800 3.3350 1.0000 ;
      RECT 2.4650 0.5700 2.5550 0.8850 ;
      RECT 2.4650 0.4800 4.6350 0.5700 ;
      RECT 2.9850 0.5700 3.0750 0.8850 ;
      RECT 3.5050 0.5700 3.5950 0.9050 ;
      RECT 4.0250 0.5700 4.1150 0.8850 ;
      RECT 4.5450 0.5700 4.6350 0.8850 ;
      RECT 4.6500 1.0950 5.5550 1.1500 ;
      RECT 3.7650 1.0500 5.5550 1.0950 ;
      RECT 0.3650 1.5850 0.4550 1.9350 ;
      RECT 0.8850 1.5850 0.9750 1.9350 ;
      RECT 1.4050 1.5850 1.4950 1.9350 ;
      RECT 1.9250 1.5850 2.0150 1.9350 ;
      RECT 2.7250 1.5850 2.8150 1.9350 ;
      RECT 3.2450 1.5850 3.3350 1.9350 ;
      RECT 3.7650 1.5850 3.8550 1.9350 ;
      RECT 3.7650 0.6800 3.8550 1.0050 ;
      RECT 4.2850 1.5850 4.3750 1.9350 ;
      RECT 4.2850 0.7500 4.3750 1.0050 ;
      RECT 0.3650 1.4950 4.7400 1.5850 ;
      RECT 4.6500 1.1500 4.7400 1.4950 ;
      RECT 3.7650 1.0050 4.7400 1.0500 ;
  END
END AND4_X4M_A12TH

MACRO AND4_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 7.8450 0.3200 ;
        RECT 0.3600 0.3200 0.4600 0.6300 ;
        RECT 0.8800 0.3200 0.9800 0.6300 ;
        RECT 1.4000 0.3200 1.5000 0.6300 ;
        RECT 5.9700 0.3200 6.0700 0.6350 ;
        RECT 6.4900 0.3200 6.5900 0.6350 ;
        RECT 7.0100 0.3200 7.1100 0.6350 ;
        RECT 7.5300 0.3200 7.6300 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 7.8450 2.7200 ;
        RECT 5.9750 1.7700 6.0650 2.0800 ;
        RECT 6.4950 1.7700 6.5850 2.0800 ;
        RECT 7.0150 1.7700 7.1050 2.0800 ;
        RECT 7.5350 1.7700 7.6250 2.0800 ;
        RECT 0.8800 1.6750 0.9800 2.0800 ;
        RECT 1.4000 1.6750 1.5000 2.0800 ;
        RECT 1.9200 1.6750 2.0200 2.0800 ;
        RECT 2.4400 1.6750 2.5400 2.0800 ;
        RECT 2.9600 1.6750 3.0600 2.0800 ;
        RECT 3.4800 1.6750 3.5800 2.0800 ;
        RECT 4.0000 1.6750 4.1000 2.0800 ;
        RECT 4.5200 1.6750 4.6200 2.0800 ;
        RECT 5.0400 1.6750 5.1400 2.0800 ;
        RECT 5.5600 1.6750 5.6600 2.0800 ;
        RECT 0.3600 1.6400 0.4600 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2500 0.9050 7.3500 1.3050 ;
        RECT 6.2300 1.3050 7.3500 1.3250 ;
        RECT 6.2300 0.8900 7.3500 0.9050 ;
        RECT 6.2300 1.3250 7.3700 1.4050 ;
        RECT 6.2300 0.8050 7.3700 0.8900 ;
        RECT 6.2300 1.4050 6.3300 1.7200 ;
        RECT 6.7500 1.4050 6.8500 1.7350 ;
        RECT 7.2700 1.4050 7.3700 1.7350 ;
        RECT 6.2300 0.4750 6.3300 0.8050 ;
        RECT 6.7500 0.4750 6.8500 0.8050 ;
        RECT 7.2700 0.4750 7.3700 0.8050 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8850 1.2500 2.3000 1.3050 ;
        RECT 1.8850 1.3050 2.9000 1.4050 ;
    END
    ANTENNAGATEAREA 0.45 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3000 1.2500 3.7000 1.3050 ;
        RECT 3.1100 1.3050 4.1600 1.4050 ;
    END
    ANTENNAGATEAREA 0.45 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4350 1.2500 4.9000 1.3050 ;
        RECT 4.4350 1.3050 5.5050 1.4050 ;
    END
    ANTENNAGATEAREA 0.45 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.2500 1.1000 1.3050 ;
        RECT 0.5250 1.3050 1.5600 1.4050 ;
    END
    ANTENNAGATEAREA 0.45 ;
  END D
  OBS
    LAYER M1 ;
      RECT 6.0500 1.1000 7.1050 1.1500 ;
      RECT 4.5250 1.0600 7.1050 1.1000 ;
      RECT 3.2250 1.5850 3.3150 1.9750 ;
      RECT 3.7450 1.5850 3.8350 1.9750 ;
      RECT 4.2650 1.5850 4.3550 1.9750 ;
      RECT 4.7850 1.5850 4.8750 1.9750 ;
      RECT 4.5250 0.6600 4.6150 1.0100 ;
      RECT 5.3050 1.5850 5.3950 1.9750 ;
      RECT 5.0450 0.6600 5.1350 1.0100 ;
      RECT 5.5600 0.4650 5.6600 1.0100 ;
      RECT 0.6250 1.4950 6.1400 1.5850 ;
      RECT 6.0500 1.1550 6.1400 1.4950 ;
      RECT 4.5250 1.0100 6.1400 1.0550 ;
      RECT 6.0500 1.1500 6.2800 1.1550 ;
      RECT 4.5250 1.0550 6.2800 1.0600 ;
      RECT 2.1850 1.5850 2.2750 1.9750 ;
      RECT 2.7050 1.5850 2.7950 1.9750 ;
      RECT 0.6250 1.5850 0.7150 1.9750 ;
      RECT 1.1450 1.5850 1.2350 1.9750 ;
      RECT 1.6650 1.5850 1.7550 1.9750 ;
      RECT 0.6250 0.8600 1.7550 0.9500 ;
      RECT 1.6650 0.5700 1.7550 0.8600 ;
      RECT 1.6650 0.4800 2.7950 0.5700 ;
      RECT 2.1850 0.5700 2.2750 0.8700 ;
      RECT 2.7050 0.5700 2.7950 0.8750 ;
      RECT 0.6250 0.5300 0.7150 0.8600 ;
      RECT 1.1450 0.5300 1.2350 0.8600 ;
      RECT 1.9250 1.0000 3.0600 1.0900 ;
      RECT 1.9250 0.6600 2.0150 1.0000 ;
      RECT 2.4450 0.6600 2.5350 1.0000 ;
      RECT 2.9650 0.6600 3.0600 1.0000 ;
      RECT 2.9700 0.5700 3.0600 0.6600 ;
      RECT 2.9700 0.4800 4.0950 0.5700 ;
      RECT 3.4850 0.5700 3.5750 0.8750 ;
      RECT 4.0050 0.5700 4.0950 0.8650 ;
      RECT 3.2250 1.0000 4.3450 1.0900 ;
      RECT 4.2550 0.9150 4.3450 1.0000 ;
      RECT 3.7450 0.6950 3.8350 1.0000 ;
      RECT 3.2250 0.6600 3.3150 1.0000 ;
      RECT 4.2550 0.5700 4.3550 0.9150 ;
      RECT 4.2550 0.4800 5.3950 0.5700 ;
      RECT 4.7850 0.5700 4.8750 0.9150 ;
      RECT 5.3050 0.5700 5.3950 0.8700 ;
  END
END AND4_X6M_A12TH

MACRO AND4_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 10.4450 0.3200 ;
        RECT 0.4400 0.3200 0.5400 0.6300 ;
        RECT 0.9600 0.3200 1.0600 0.6300 ;
        RECT 1.4800 0.3200 1.5800 0.6300 ;
        RECT 2.0000 0.3200 2.1000 0.6300 ;
        RECT 8.1300 0.3200 8.2300 0.6350 ;
        RECT 8.6500 0.3200 8.7500 0.6350 ;
        RECT 9.1700 0.3200 9.2700 0.6350 ;
        RECT 9.6900 0.3200 9.7900 0.6350 ;
        RECT 10.2100 0.3200 10.3100 0.6350 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 10.4450 2.7200 ;
        RECT 8.1350 1.7700 8.2250 2.0800 ;
        RECT 8.6550 1.7700 8.7450 2.0800 ;
        RECT 9.1750 1.7700 9.2650 2.0800 ;
        RECT 9.6950 1.7700 9.7850 2.0800 ;
        RECT 10.2150 1.7700 10.3050 2.0800 ;
        RECT 0.9600 1.6750 1.0600 2.0800 ;
        RECT 1.4800 1.6750 1.5800 2.0800 ;
        RECT 2.0000 1.6750 2.1000 2.0800 ;
        RECT 2.5200 1.6750 2.6200 2.0800 ;
        RECT 3.0400 1.6750 3.1400 2.0800 ;
        RECT 3.5600 1.6750 3.6600 2.0800 ;
        RECT 4.0800 1.6750 4.1800 2.0800 ;
        RECT 4.6000 1.6750 4.7000 2.0800 ;
        RECT 5.1200 1.6750 5.2200 2.0800 ;
        RECT 5.6400 1.6750 5.7400 2.0800 ;
        RECT 6.1600 1.6750 6.2600 2.0800 ;
        RECT 6.6800 1.6750 6.7800 2.0800 ;
        RECT 7.2000 1.6750 7.3000 2.0800 ;
        RECT 7.7200 1.6750 7.8200 2.0800 ;
        RECT 0.4400 1.6400 0.5400 2.0800 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3000 1.2500 1.7000 1.3050 ;
        RECT 0.9000 1.3050 1.9000 1.4050 ;
    END
    ANTENNAGATEAREA 0.609 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.3000 1.2500 6.7000 1.3050 ;
        RECT 6.3000 1.3050 7.3400 1.4050 ;
    END
    ANTENNAGATEAREA 0.609 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9000 1.2500 5.3000 1.3050 ;
        RECT 4.5000 1.3050 5.5300 1.4050 ;
    END
    ANTENNAGATEAREA 0.609 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7000 1.2500 3.1000 1.3050 ;
        RECT 2.7000 1.3050 3.7050 1.4050 ;
    END
    ANTENNAGATEAREA 0.609 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.4350 1.4200 9.5650 1.7350 ;
        RECT 8.3750 1.2900 10.0650 1.4200 ;
        RECT 8.3750 1.4200 8.5050 1.7200 ;
        RECT 8.8950 1.4200 9.0250 1.7350 ;
        RECT 9.9350 1.4200 10.0650 1.7350 ;
        RECT 9.9350 0.9200 10.0650 1.2900 ;
        RECT 8.3750 0.7900 10.0650 0.9200 ;
        RECT 8.3750 0.4750 8.5050 0.7900 ;
        RECT 8.8950 0.4750 9.0250 0.7900 ;
        RECT 9.4150 0.4750 9.5450 0.7900 ;
        RECT 9.9350 0.4750 10.0650 0.7900 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.7050 0.8600 2.3550 0.9500 ;
      RECT 2.2650 0.5700 2.3550 0.8600 ;
      RECT 2.2650 0.4800 3.9150 0.5700 ;
      RECT 2.7850 0.5700 2.8750 0.9100 ;
      RECT 3.3050 0.5700 3.3950 0.9100 ;
      RECT 3.8250 0.5700 3.9150 0.8750 ;
      RECT 0.7050 0.5300 0.7950 0.8600 ;
      RECT 1.2250 0.5500 1.3150 0.8600 ;
      RECT 1.7450 0.5300 1.8350 0.8600 ;
      RECT 2.5250 1.0000 4.1750 1.0900 ;
      RECT 2.5250 0.6600 2.6150 1.0000 ;
      RECT 3.0450 0.6600 3.1350 1.0000 ;
      RECT 3.5650 0.6600 3.6550 1.0000 ;
      RECT 4.0850 0.5700 4.1750 1.0000 ;
      RECT 4.0850 0.4800 5.7350 0.5700 ;
      RECT 4.6050 0.5700 4.6950 0.8700 ;
      RECT 5.1250 0.5700 5.2150 0.8750 ;
      RECT 5.6450 0.5700 5.7350 0.8650 ;
      RECT 4.3450 1.0000 5.9850 1.0900 ;
      RECT 5.8950 0.9150 5.9850 1.0000 ;
      RECT 5.3850 0.6950 5.4750 1.0000 ;
      RECT 4.8650 0.6750 4.9550 1.0000 ;
      RECT 4.3450 0.6600 4.4350 1.0000 ;
      RECT 5.8950 0.5700 5.9950 0.9150 ;
      RECT 5.8950 0.4800 7.5550 0.5700 ;
      RECT 6.4250 0.5700 6.5150 0.9150 ;
      RECT 6.9450 0.5700 7.0350 0.8700 ;
      RECT 7.4650 0.5700 7.5550 0.8700 ;
      RECT 8.1750 1.1000 9.2650 1.1550 ;
      RECT 6.1650 1.0550 9.2650 1.1000 ;
      RECT 6.4250 1.5850 6.5150 1.9750 ;
      RECT 6.9450 1.5850 7.0350 1.9750 ;
      RECT 6.6800 0.6900 6.7800 1.0100 ;
      RECT 7.4650 1.5850 7.5550 1.9750 ;
      RECT 7.2000 0.6600 7.3000 1.0100 ;
      RECT 7.7200 0.4650 7.8200 1.0100 ;
      RECT 0.7050 1.4950 8.2650 1.5850 ;
      RECT 8.1750 1.1550 8.2650 1.4950 ;
      RECT 6.1650 1.0100 8.2650 1.0550 ;
      RECT 4.8650 1.5850 4.9550 1.9750 ;
      RECT 5.3850 1.5850 5.4750 1.9750 ;
      RECT 5.9050 1.5850 5.9950 1.9750 ;
      RECT 6.1650 0.6600 6.2550 1.0100 ;
      RECT 2.7850 1.5850 2.8750 1.9750 ;
      RECT 3.3050 1.5850 3.3950 1.9750 ;
      RECT 3.8250 1.5850 3.9150 1.9750 ;
      RECT 4.3450 1.5850 4.4350 1.9750 ;
      RECT 1.2250 1.5850 1.3150 1.9550 ;
      RECT 1.7450 1.5850 1.8350 1.9550 ;
      RECT 2.2650 1.5850 2.3550 1.9550 ;
      RECT 0.7050 1.5850 0.7950 1.9750 ;
  END
END AND4_X8M_A12TH

MACRO ANTENNA2_A12TH
  CLASS CORE ANTENNACELL ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 0.4450 0.3200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 0.4450 2.7200 ;
    END
  END VDD

  PIN A
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.0600 0.6100 0.3500 0.7900 ;
    END
    ANTENNADIFFAREA 0.06 ;
  END A
END ANTENNA2_A12TH

MACRO AO1B2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6450 0.3200 0.7350 0.6950 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1800 1.7050 1.2700 2.0800 ;
        RECT 0.1250 1.6700 0.2150 2.0800 ;
        RECT 0.6450 1.6700 0.7350 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7700 0.5500 1.1900 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8450 0.7850 0.9550 1.1800 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END A0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6450 1.3500 1.5000 ;
        RECT 0.9500 1.5000 1.3500 1.6000 ;
        RECT 1.1200 0.5550 1.3500 0.6450 ;
        RECT 0.9500 1.6000 1.0500 1.6900 ;
        RECT 0.8800 1.6900 1.0500 1.9800 ;
    END
    ANTENNADIFFAREA 0.162925 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2550 1.3000 1.1550 1.3900 ;
      RECT 0.3850 1.3900 0.4750 1.8850 ;
      RECT 0.2550 0.6500 0.3450 1.3000 ;
      RECT 0.0650 0.5600 0.3450 0.6500 ;
  END
END AO1B2_X0P5M_A12TH

MACRO AO1B2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6450 0.3200 0.7350 0.7150 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1800 1.7500 1.2700 2.0800 ;
        RECT 0.1200 1.6800 0.2200 2.0800 ;
        RECT 0.6450 1.6350 0.7350 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0550 0.1600 1.4550 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.8050 0.5550 1.1900 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8450 0.8050 0.9550 1.1900 ;
    END
    ANTENNAGATEAREA 0.0684 ;
  END A0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.7500 1.3500 1.5300 ;
        RECT 0.9150 1.5300 1.3500 1.6300 ;
        RECT 1.1400 0.4600 1.3500 0.7500 ;
        RECT 0.9150 1.6300 1.0150 1.9600 ;
    END
    ANTENNADIFFAREA 0.230725 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2550 1.3200 1.1450 1.4100 ;
      RECT 0.3850 1.4100 0.4750 1.7950 ;
      RECT 0.2550 0.7000 0.3450 1.3200 ;
      RECT 0.0650 0.6100 0.3450 0.7000 ;
  END
END AO1B2_X0P7M_A12TH

MACRO AO1B2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6350 0.3200 0.7350 0.6300 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9850 0.1600 1.4000 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.7700 0.5500 1.2300 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7350 0.8500 1.0400 0.9500 ;
        RECT 0.7350 0.9500 0.8350 1.2300 ;
    END
    ANTENNAGATEAREA 0.0969 ;
  END A0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9700 1.3500 1.5500 ;
        RECT 0.8950 1.5500 1.3500 1.6500 ;
        RECT 1.1550 0.8700 1.3500 0.9700 ;
        RECT 0.8950 1.6500 0.9950 1.9600 ;
        RECT 1.1550 0.5400 1.2550 0.8700 ;
    END
    ANTENNADIFFAREA 0.32685 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6350 1.7500 0.7350 2.0800 ;
        RECT 1.1550 1.7500 1.2550 2.0800 ;
        RECT 0.0900 1.5100 0.1900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2550 1.3400 1.0750 1.4300 ;
      RECT 0.9850 1.0700 1.0750 1.3400 ;
      RECT 0.3550 1.4300 0.4450 1.9200 ;
      RECT 0.2550 0.8650 0.3450 1.3400 ;
      RECT 0.0900 0.7750 0.3450 0.8650 ;
      RECT 0.0900 0.6550 0.1900 0.7750 ;
  END
END AO1B2_X1M_A12TH

MACRO AO1B2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.6800 0.3200 0.7700 0.7500 ;
        RECT 1.7500 0.3200 1.8400 0.6750 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.2150 1.7600 1.3050 2.0800 ;
        RECT 1.7500 1.7600 1.8400 2.0800 ;
        RECT 0.1600 1.6800 0.2500 2.0800 ;
        RECT 0.6800 1.6150 0.7700 2.0800 ;
    END
  END VDD

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1600 1.5000 ;
    END
    ANTENNAGATEAREA 0.0564 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8950 0.5900 1.1950 ;
    END
    ANTENNAGATEAREA 0.0564 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8800 1.0500 1.7500 1.1500 ;
        RECT 1.6450 1.1500 1.7500 1.4200 ;
        RECT 0.8800 0.9400 0.9800 1.0500 ;
    END
    ANTENNAGATEAREA 0.1368 ;
  END A0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8950 1.9500 1.5400 ;
        RECT 0.9550 1.5400 1.9500 1.6400 ;
        RECT 1.2100 0.7950 1.9500 0.8950 ;
        RECT 0.9550 1.6400 1.0450 1.9550 ;
        RECT 1.4900 1.6400 1.5800 1.9550 ;
        RECT 1.2100 0.4400 1.3100 0.7950 ;
    END
    ANTENNADIFFAREA 0.355175 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2550 1.3150 1.4700 1.4050 ;
      RECT 0.4200 1.4050 0.5100 1.9600 ;
      RECT 0.2550 0.7000 0.3450 1.3150 ;
      RECT 0.1200 0.6100 0.3450 0.7000 ;
      RECT 0.1200 0.4100 0.2900 0.6100 ;
  END
END AO1B2_X1P4M_A12TH

MACRO AO1B2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.2000 1.7950 1.2900 2.0800 ;
        RECT 1.7350 1.7950 1.8250 2.0800 ;
        RECT 0.1450 1.7550 0.2350 2.0800 ;
        RECT 0.6650 1.7550 0.7550 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.6250 0.3200 0.7950 0.5100 ;
        RECT 1.6950 0.3200 1.8650 0.5300 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0900 0.1600 1.5100 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B0

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9700 0.5700 1.3900 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8500 1.7500 0.9500 ;
        RECT 0.8500 0.9500 0.9500 1.2600 ;
        RECT 1.6500 0.9500 1.7500 1.2600 ;
    END
    ANTENNAGATEAREA 0.1938 ;
  END A0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.7500 1.9500 1.5700 ;
        RECT 0.9350 1.5700 1.9500 1.6700 ;
        RECT 1.1650 0.6500 1.9500 0.7500 ;
        RECT 0.9350 1.6700 1.0350 1.9600 ;
        RECT 1.4750 1.6700 1.5650 1.9600 ;
        RECT 1.1650 0.4600 1.3350 0.6500 ;
    END
    ANTENNADIFFAREA 0.50355 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.0700 1.1100 1.4750 1.2000 ;
      RECT 0.4050 1.5250 0.7500 1.6150 ;
      RECT 0.6600 1.4600 0.7500 1.5250 ;
      RECT 0.6600 0.7200 0.7500 1.3700 ;
      RECT 0.1000 0.6300 0.7500 0.7200 ;
      RECT 0.6600 1.3700 1.1600 1.4600 ;
      RECT 1.0700 1.2000 1.1600 1.3700 ;
      RECT 0.4050 1.6150 0.4950 1.9600 ;
      RECT 0.1000 0.4300 0.2700 0.6300 ;
  END
END AO1B2_X2M_A12TH

MACRO AO1B2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.1400 0.3200 0.2300 0.6300 ;
        RECT 1.1400 0.3200 1.3100 0.5300 ;
        RECT 2.2100 0.3200 2.3800 0.5300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 1.7150 1.7950 1.8050 2.0800 ;
        RECT 2.2500 1.7950 2.3400 2.0800 ;
        RECT 2.7700 1.7950 2.8600 2.0800 ;
        RECT 0.1400 1.7550 0.2300 2.0800 ;
        RECT 0.6600 1.7550 0.7500 2.0800 ;
        RECT 1.1800 1.7550 1.2700 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1550 0.8500 1.1000 0.9500 ;
        RECT 1.0000 0.9500 1.1000 1.3700 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3800 0.8500 2.2150 0.9500 ;
        RECT 2.1150 0.9500 2.2150 1.0500 ;
        RECT 1.3800 0.9500 1.4800 1.2500 ;
        RECT 2.1150 1.0500 2.5250 1.1500 ;
    END
    ANTENNAGATEAREA 0.2907 ;
  END A0N

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4700 1.2500 0.8900 1.3500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8500 0.7500 2.9500 1.5700 ;
        RECT 1.4500 1.5700 2.9500 1.6700 ;
        RECT 1.6800 0.6500 2.9500 0.7500 ;
        RECT 1.4500 1.6700 1.5500 1.9600 ;
        RECT 1.9900 1.6700 2.0800 1.9600 ;
        RECT 2.5100 1.6700 2.6000 1.9600 ;
        RECT 1.6800 0.4600 1.8500 0.6500 ;
        RECT 2.7300 0.4600 2.9000 0.6500 ;
    END
    ANTENNADIFFAREA 0.8304 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.1950 1.3600 2.7550 1.4500 ;
      RECT 2.6650 1.0500 2.7550 1.3600 ;
      RECT 0.4000 1.6300 0.4900 1.9100 ;
      RECT 0.9200 1.6300 1.0100 1.9100 ;
      RECT 0.6600 0.4750 0.7500 0.6550 ;
      RECT 0.4000 1.5400 1.2850 1.6300 ;
      RECT 1.1950 1.4500 1.2850 1.5400 ;
      RECT 1.1950 0.7450 1.2850 1.3600 ;
      RECT 0.6600 0.6550 1.2850 0.7450 ;
      RECT 1.8950 1.2000 1.9850 1.3600 ;
      RECT 1.5950 1.1100 1.9850 1.2000 ;
  END
END AO1B2_X3M_A12TH

MACRO AO1B2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6300 ;
        RECT 1.0800 0.3200 1.2500 0.5500 ;
        RECT 2.1500 0.3200 2.3200 0.5300 ;
        RECT 3.2250 0.3200 3.3250 0.4450 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.6550 1.7900 1.7450 2.0800 ;
        RECT 2.1900 1.7900 2.2800 2.0800 ;
        RECT 2.7100 1.7900 2.8000 2.0800 ;
        RECT 3.2300 1.7900 3.3200 2.0800 ;
        RECT 0.0800 1.7550 0.1700 2.0800 ;
        RECT 0.6000 1.7550 0.6900 2.0800 ;
        RECT 1.1200 1.7550 1.2100 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 0.8500 1.0300 0.9500 ;
        RECT 0.2550 0.9500 0.3550 1.1200 ;
        RECT 0.9300 0.9500 1.0300 1.2800 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END B1

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3200 0.8500 3.1500 0.9500 ;
        RECT 2.0600 0.9500 2.1600 1.0500 ;
        RECT 1.3200 0.9500 1.4200 1.2600 ;
        RECT 3.0500 0.9500 3.1500 1.2600 ;
        RECT 2.0600 1.0500 2.4500 1.1500 ;
    END
    ANTENNAGATEAREA 0.3876 ;
  END A0N

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.2500 0.8300 1.3500 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END B0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 0.7500 3.3500 1.5700 ;
        RECT 1.3900 1.5700 3.3500 1.6700 ;
        RECT 1.6200 0.6500 3.3500 0.7500 ;
        RECT 1.3900 1.6700 1.4900 1.9600 ;
        RECT 1.9300 1.6700 2.0200 1.9600 ;
        RECT 2.4500 1.6700 2.5400 1.9600 ;
        RECT 2.9700 1.6700 3.0600 1.9600 ;
        RECT 1.6200 0.4600 1.7900 0.6500 ;
        RECT 2.6700 0.4550 2.8400 0.6500 ;
    END
    ANTENNADIFFAREA 0.99555 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 2.5700 1.1100 2.9450 1.2000 ;
      RECT 1.1200 1.3600 2.6600 1.4500 ;
      RECT 2.5700 1.2000 2.6600 1.3600 ;
      RECT 0.8600 1.6150 0.9500 1.9600 ;
      RECT 0.3400 1.5250 1.2100 1.6150 ;
      RECT 1.1200 1.4500 1.2100 1.5250 ;
      RECT 1.1200 0.7450 1.2100 1.3600 ;
      RECT 0.5600 0.6550 1.2100 0.7450 ;
      RECT 1.5300 1.2000 1.6200 1.3600 ;
      RECT 1.5300 1.1100 1.9200 1.2000 ;
      RECT 0.3400 1.6150 0.4300 1.9600 ;
      RECT 0.5600 0.4550 0.7300 0.6550 ;
  END
END AO1B2_X4M_A12TH

MACRO AO1B2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.6200 0.3200 0.7100 0.7100 ;
        RECT 1.6600 0.3200 1.7500 0.7100 ;
        RECT 2.7300 0.3200 2.8200 0.5600 ;
        RECT 3.7700 0.3200 3.8600 0.5600 ;
        RECT 4.8100 0.3200 4.9000 0.5600 ;
    END
  END VSS

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1150 1.0500 1.3500 1.1500 ;
    END
    ANTENNAGATEAREA 0.2304 ;
  END B0

  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8550 0.8500 4.7500 0.9500 ;
        RECT 2.5950 0.9500 2.6950 1.0600 ;
        RECT 1.8550 0.9500 1.9550 1.2600 ;
        RECT 3.6350 0.9500 3.7350 1.0600 ;
        RECT 4.6500 0.9500 4.7500 1.2600 ;
        RECT 2.5950 1.0600 2.9850 1.1600 ;
        RECT 3.6350 1.0600 4.0250 1.1600 ;
    END
    ANTENNAGATEAREA 0.5814 ;
  END A0N

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 2.1950 1.7900 2.2850 2.0800 ;
        RECT 2.7300 1.7900 2.8200 2.0800 ;
        RECT 3.2500 1.7900 3.3400 2.0800 ;
        RECT 3.7700 1.7900 3.8600 2.0800 ;
        RECT 4.2900 1.7900 4.3800 2.0800 ;
        RECT 4.8100 1.7900 4.9000 2.0800 ;
        RECT 0.1000 1.7550 0.1900 2.0800 ;
        RECT 0.6200 1.7550 0.7100 2.0800 ;
        RECT 1.1400 1.7550 1.2300 2.0800 ;
        RECT 1.6600 1.7550 1.7500 2.0800 ;
    END
  END VDD

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.1400 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2304 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.7500 4.9500 1.5700 ;
        RECT 1.9300 1.5700 4.9500 1.6700 ;
        RECT 2.1600 0.6500 4.9500 0.7500 ;
        RECT 1.9300 1.6700 2.0300 1.9600 ;
        RECT 2.4700 1.6700 2.5600 1.9600 ;
        RECT 2.9900 1.6700 3.0800 1.9600 ;
        RECT 3.5100 1.6700 3.6000 1.9600 ;
        RECT 4.0300 1.6700 4.1200 1.9600 ;
        RECT 4.5500 1.6700 4.6400 1.9600 ;
        RECT 2.1600 0.4600 2.3300 0.6500 ;
        RECT 3.2100 0.4600 3.3800 0.6500 ;
        RECT 4.2500 0.4600 4.4200 0.6500 ;
    END
    ANTENNADIFFAREA 1.48755 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 4.1450 1.1100 4.5300 1.2000 ;
      RECT 1.6550 1.3600 4.2350 1.4500 ;
      RECT 4.1450 1.2000 4.2350 1.3600 ;
      RECT 0.1000 0.4700 0.1900 0.8100 ;
      RECT 0.3600 1.6250 0.4500 1.9550 ;
      RECT 0.8800 1.6250 0.9700 1.9550 ;
      RECT 1.4000 1.6250 1.4900 1.9550 ;
      RECT 1.1400 0.4700 1.2300 0.8100 ;
      RECT 0.3600 1.5350 1.7450 1.6250 ;
      RECT 1.6550 1.4500 1.7450 1.5350 ;
      RECT 1.6550 0.9000 1.7450 1.3600 ;
      RECT 0.1000 0.8100 1.7450 0.9000 ;
      RECT 2.0700 1.2000 2.1600 1.3600 ;
      RECT 2.0700 1.1100 2.4600 1.2000 ;
      RECT 3.1050 1.2000 3.1950 1.3600 ;
      RECT 3.1050 1.1100 3.5050 1.2000 ;
  END
END AO1B2_X6M_A12TH

MACRO AO21B_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6450 0.3200 0.7350 0.6950 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.6300 1.3500 1.5000 ;
        RECT 0.9150 1.5000 1.3500 1.6000 ;
        RECT 1.1200 0.5400 1.3500 0.6300 ;
        RECT 0.9150 1.6000 1.0150 1.9900 ;
    END
    ANTENNADIFFAREA 0.162925 ;
  END Y

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0200 0.9750 1.1500 1.3450 ;
    END
    ANTENNAGATEAREA 0.0483 ;
  END B0N

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.3800 0.7500 1.5850 ;
        RECT 0.4500 1.2800 0.7500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0550 0.1600 1.4500 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.6050 1.6900 0.7750 2.0800 ;
        RECT 1.1800 1.6900 1.2700 2.0800 ;
        RECT 0.1150 1.6750 0.2250 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2550 0.8300 0.9100 0.9200 ;
      RECT 0.2550 0.9200 0.3450 1.5000 ;
      RECT 0.2550 0.6350 0.3450 0.8300 ;
      RECT 0.0650 0.5450 0.3450 0.6350 ;
      RECT 0.3850 1.5900 0.4750 1.8400 ;
      RECT 0.2550 1.5000 0.4750 1.5900 ;
  END
END AO21B_X0P5M_A12TH

MACRO AO21B_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6450 0.3200 0.7350 0.7200 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.0850 1.8150 0.1750 2.0800 ;
        RECT 1.1800 1.7500 1.2700 2.0800 ;
        RECT 0.6450 1.6800 0.7350 2.0800 ;
        RECT 0.0850 1.7250 0.2750 1.8150 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0800 0.1600 1.5150 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 1.3500 0.7500 1.5900 ;
        RECT 0.4700 1.2500 0.7500 1.3500 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0200 0.9850 1.1500 1.3850 ;
    END
    ANTENNAGATEAREA 0.0684 ;
  END B0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.8100 1.3500 1.5200 ;
        RECT 0.9150 1.5200 1.3500 1.6200 ;
        RECT 1.1800 0.4400 1.3500 0.8100 ;
        RECT 0.9150 1.6200 1.0150 1.9800 ;
    END
    ANTENNADIFFAREA 0.230725 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2550 0.8100 0.8400 0.9000 ;
      RECT 0.7500 0.9000 0.8400 1.1000 ;
      RECT 0.2550 0.9000 0.3450 1.4950 ;
      RECT 0.2550 0.7000 0.3450 0.8100 ;
      RECT 0.0650 0.6100 0.3450 0.7000 ;
      RECT 0.3850 1.5850 0.4750 1.8250 ;
      RECT 0.2550 1.4950 0.4750 1.5850 ;
  END
END AO21B_X0P7M_A12TH

MACRO AO21B_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6450 0.3200 0.7350 0.5000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.1250 1.7800 0.2150 2.0800 ;
        RECT 0.6450 1.7800 0.7350 2.0800 ;
        RECT 1.1800 1.7750 1.2700 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2450 0.1600 1.6700 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9800 0.5600 1.3900 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2400 1.0500 1.3500 1.4350 ;
    END
    ANTENNAGATEAREA 0.0969 ;
  END B0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9300 1.1500 1.4500 ;
        RECT 0.9150 1.4500 1.1500 1.5500 ;
        RECT 1.0500 0.8300 1.2750 0.9300 ;
        RECT 0.9150 1.5500 1.0150 1.8600 ;
        RECT 1.1750 0.5200 1.2750 0.8300 ;
    END
    ANTENNADIFFAREA 0.32685 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.3850 1.5850 0.7450 1.6750 ;
      RECT 0.6550 1.2400 0.7450 1.5850 ;
      RECT 0.6550 1.0700 0.8100 1.2400 ;
      RECT 0.6550 0.7000 0.7450 1.0700 ;
      RECT 0.1250 0.6100 0.7450 0.7000 ;
      RECT 0.3850 1.6750 0.4750 1.8550 ;
      RECT 0.1250 0.4250 0.2150 0.6100 ;
  END
END AO21B_X1M_A12TH

MACRO AO21B_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.6450 0.3200 0.7350 0.7200 ;
        RECT 1.7150 0.3200 1.8050 0.6700 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 1.1800 1.7650 1.2700 2.0800 ;
        RECT 1.7150 1.7650 1.8050 2.0800 ;
        RECT 0.1250 1.6800 0.2150 2.0800 ;
        RECT 0.6450 1.6200 0.7350 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.1000 0.1600 1.5200 ;
    END
    ANTENNAGATEAREA 0.0564 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.8050 0.5600 1.1900 ;
    END
    ANTENNAGATEAREA 0.0564 ;
  END A1

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.0500 1.4600 1.1500 ;
    END
    ANTENNAGATEAREA 0.1368 ;
  END B0N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.8900 1.9500 1.5450 ;
        RECT 0.9200 1.5450 1.9500 1.6450 ;
        RECT 1.1750 0.7900 1.9500 0.8900 ;
        RECT 0.9200 1.6450 1.0200 1.9600 ;
        RECT 1.4550 1.6450 1.5450 1.9600 ;
        RECT 1.1750 0.4400 1.2750 0.7900 ;
    END
    ANTENNADIFFAREA 0.355175 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 0.2550 1.3300 1.7450 1.4200 ;
      RECT 1.6550 1.0100 1.7450 1.3300 ;
      RECT 0.3850 1.4200 0.4750 1.9600 ;
      RECT 0.2550 0.9000 0.3450 1.3300 ;
      RECT 0.1250 0.8100 0.3450 0.9000 ;
      RECT 0.1250 0.4400 0.2150 0.8100 ;
  END
END AO21B_X1P4M_A12TH

MACRO AO21B_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.6050 1.8800 0.7750 2.0800 ;
        RECT 0.1250 1.7550 0.2150 2.0800 ;
        RECT 1.1800 1.7550 1.2700 2.0800 ;
        RECT 1.7150 1.7550 1.8050 2.0800 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.6050 0.3200 0.7750 0.5250 ;
        RECT 1.6750 0.3200 1.8450 0.5300 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8500 0.7500 1.9500 1.4750 ;
        RECT 0.9150 1.4750 1.9500 1.5750 ;
        RECT 1.1450 0.6500 1.9500 0.7500 ;
        RECT 0.9150 1.5750 1.0150 1.8850 ;
        RECT 1.4550 1.5750 1.5450 1.8850 ;
        RECT 1.1450 0.4400 1.3150 0.6500 ;
    END
    ANTENNADIFFAREA 0.50355 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0800 0.5900 1.4100 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0850 0.1600 1.4700 ;
    END
    ANTENNAGATEAREA 0.0756 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0400 1.0500 1.4600 1.1500 ;
    END
    ANTENNAGATEAREA 0.1938 ;
  END B0N
  OBS
    LAYER M1 ;
      RECT 0.7200 0.8550 1.7500 0.9450 ;
      RECT 1.6600 0.9450 1.7500 1.2600 ;
      RECT 0.3450 1.7700 0.5150 1.9750 ;
      RECT 0.0850 0.4100 0.2550 0.6300 ;
      RECT 0.3450 1.6800 0.8100 1.7700 ;
      RECT 0.7200 0.9450 0.8100 1.6800 ;
      RECT 0.7200 0.7200 0.8100 0.8550 ;
      RECT 0.0850 0.6300 0.8100 0.7200 ;
  END
END AO21B_X2M_A12TH

MACRO AO21B_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6050 ;
        RECT 1.0900 0.3200 1.2600 0.5550 ;
        RECT 2.1100 0.3200 2.2000 0.6300 ;
    END
  END VSS

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4550 1.0800 1.8250 1.1800 ;
        RECT 1.6100 1.0500 1.8250 1.0800 ;
        RECT 1.7350 1.0200 1.8250 1.0500 ;
        RECT 1.7350 0.9300 2.5600 1.0200 ;
        RECT 2.4700 1.0200 2.5600 1.2400 ;
    END
    ANTENNAGATEAREA 0.2907 ;
  END B0N

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.0500 1.0400 1.1500 ;
        RECT 0.2100 0.9300 0.3100 1.0500 ;
        RECT 0.9500 0.9300 1.0400 1.0500 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4250 0.8500 0.8100 0.9600 ;
    END
    ANTENNAGATEAREA 0.1164 ;
  END A0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3300 1.4500 2.7500 1.5500 ;
        RECT 1.3300 1.5500 1.4200 1.8800 ;
        RECT 1.8500 1.5500 1.9400 1.8800 ;
        RECT 2.3700 1.5500 2.4600 1.8800 ;
        RECT 2.6500 0.8400 2.7500 1.4500 ;
        RECT 1.5900 0.7500 2.7500 0.8400 ;
        RECT 1.5900 0.4500 1.6800 0.7500 ;
        RECT 2.6300 0.4500 2.7200 0.7500 ;
    END
    ANTENNADIFFAREA 0.7842 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 0.0950 1.9900 0.1850 2.0800 ;
        RECT 0.9950 1.9900 1.0850 2.0800 ;
        RECT 1.5900 1.7350 1.6800 2.0800 ;
        RECT 2.1100 1.7350 2.2000 2.0800 ;
        RECT 2.6300 1.7350 2.7200 2.0800 ;
        RECT 0.5850 1.4450 0.6750 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3250 1.2650 1.3350 1.2700 ;
      RECT 0.3250 1.2700 2.0050 1.3550 ;
      RECT 0.3250 1.3550 0.4150 1.7500 ;
      RECT 0.5450 0.6700 1.2200 0.7600 ;
      RECT 0.5450 0.4250 0.7150 0.6700 ;
      RECT 0.8450 1.3550 0.9350 1.7500 ;
      RECT 1.1300 1.3550 2.0050 1.3600 ;
      RECT 1.1300 0.7600 1.2200 1.0500 ;
      RECT 1.9150 1.2000 2.0050 1.2700 ;
      RECT 1.9150 1.1100 2.3350 1.2000 ;
      RECT 1.1300 1.0500 1.3350 1.3600 ;
  END
END AO21B_X3M_A12TH

MACRO AO21B_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7050 ;
        RECT 1.1500 0.3200 1.2400 0.7250 ;
        RECT 2.1900 0.3200 2.2800 0.5600 ;
        RECT 3.2300 0.3200 3.3200 0.5600 ;
    END
  END VSS

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 1.0500 0.7950 1.1600 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5200 1.0500 1.8950 1.1800 ;
        RECT 1.8050 0.9500 1.8950 1.0500 ;
        RECT 1.8050 0.8500 2.5950 0.9500 ;
        RECT 2.5050 0.9500 2.5950 1.0900 ;
        RECT 2.5050 1.0900 2.9350 1.1800 ;
    END
    ANTENNAGATEAREA 0.3876 ;
  END B0N

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2100 1.2500 1.0150 1.3500 ;
        RECT 0.2100 1.2350 0.3000 1.2500 ;
        RECT 0.9250 1.2350 1.0150 1.2500 ;
        RECT 0.0900 1.1450 0.3000 1.2350 ;
        RECT 0.9250 1.1450 1.1350 1.2350 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.4500 3.3500 1.5500 ;
        RECT 1.4100 1.5500 1.5000 1.8800 ;
        RECT 1.9300 1.5500 2.0200 1.8800 ;
        RECT 2.4500 1.5500 2.5400 1.8800 ;
        RECT 2.9700 1.5500 3.0600 1.8800 ;
        RECT 3.2500 0.7500 3.3500 1.4500 ;
        RECT 1.6300 0.6550 3.3500 0.7500 ;
        RECT 1.6300 0.6500 2.8400 0.6550 ;
        RECT 1.6300 0.4100 1.8000 0.6500 ;
        RECT 2.6700 0.4100 2.8400 0.6500 ;
    END
    ANTENNADIFFAREA 0.984 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 1.6700 1.7500 1.7600 2.0800 ;
        RECT 2.1900 1.7500 2.2800 2.0800 ;
        RECT 2.7100 1.7500 2.8000 2.0800 ;
        RECT 3.2300 1.7500 3.3200 2.0800 ;
        RECT 0.6000 1.6200 0.6900 2.0800 ;
        RECT 1.1500 1.6200 1.2400 2.0800 ;
        RECT 0.0800 1.5500 0.1700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.3250 1.2700 3.1600 1.3600 ;
      RECT 3.0700 1.0500 3.1600 1.2700 ;
      RECT 2.0450 1.1100 2.4150 1.2000 ;
      RECT 2.3250 1.2000 2.4150 1.2700 ;
      RECT 0.3400 1.5300 0.4300 1.8700 ;
      RECT 0.8600 1.5300 0.9500 1.8700 ;
      RECT 0.6000 0.4950 0.6900 0.8650 ;
      RECT 0.3400 1.4400 1.3200 1.5300 ;
      RECT 1.2300 1.3600 1.3200 1.4400 ;
      RECT 1.2300 1.0500 1.3550 1.2700 ;
      RECT 1.2300 0.9550 1.3200 1.0500 ;
      RECT 0.6000 0.8650 1.3200 0.9550 ;
      RECT 1.2300 1.2700 2.1350 1.3600 ;
      RECT 2.0450 1.2000 2.1350 1.2700 ;
  END
END AO21B_X4M_A12TH

MACRO AO21B_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.6200 0.3200 0.7100 0.6900 ;
        RECT 1.6600 0.3200 1.7500 0.6900 ;
        RECT 2.7300 0.3200 2.8200 0.5600 ;
        RECT 3.7700 0.3200 3.8600 0.5600 ;
        RECT 4.8100 0.3200 4.9000 0.5600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.1000 1.7550 0.1900 2.0800 ;
        RECT 0.6200 1.7550 0.7100 2.0800 ;
        RECT 1.1400 1.7550 1.2300 2.0800 ;
        RECT 1.6600 1.7550 1.7500 2.0800 ;
        RECT 2.1950 1.7550 2.2850 2.0800 ;
        RECT 2.7300 1.7550 2.8200 2.0800 ;
        RECT 3.2500 1.7550 3.3400 2.0800 ;
        RECT 3.7700 1.7550 3.8600 2.0800 ;
        RECT 4.2900 1.7550 4.3800 2.0800 ;
        RECT 4.8100 1.7550 4.9000 2.0800 ;
    END
  END VDD

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1150 1.0500 1.3500 1.1500 ;
    END
    ANTENNAGATEAREA 0.2304 ;
  END A0

  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3200 0.8500 4.2150 0.9500 ;
        RECT 2.3200 0.9500 2.4200 1.0500 ;
        RECT 3.3750 0.9500 3.4750 1.0500 ;
        RECT 4.1150 0.9500 4.2150 1.0500 ;
        RECT 2.0100 1.0500 2.4200 1.1500 ;
        RECT 3.0700 1.0500 3.4750 1.1500 ;
        RECT 4.1150 1.0500 4.5150 1.1500 ;
    END
    ANTENNAGATEAREA 0.5814 ;
  END B0N

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.2500 1.5800 1.3500 ;
        RECT 1.4750 1.1400 1.5800 1.2500 ;
    END
    ANTENNAGATEAREA 0.2304 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.7500 4.9500 1.4500 ;
        RECT 1.9300 1.4500 4.9500 1.5500 ;
        RECT 2.1600 0.6500 4.9500 0.7500 ;
        RECT 1.9300 1.5500 2.0300 1.8800 ;
        RECT 2.4700 1.5500 2.5600 1.8800 ;
        RECT 2.9900 1.5500 3.0800 1.8800 ;
        RECT 3.5100 1.5500 3.6000 1.8800 ;
        RECT 4.0300 1.5500 4.1200 1.8800 ;
        RECT 4.5500 1.5500 4.6400 1.8800 ;
        RECT 2.1600 0.4550 2.3300 0.6500 ;
        RECT 3.2100 0.4550 3.3800 0.6500 ;
        RECT 4.2500 0.4550 4.4200 0.6500 ;
    END
    ANTENNADIFFAREA 1.48755 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.7350 1.2500 4.7500 1.3500 ;
      RECT 4.6500 1.0500 4.7500 1.2500 ;
      RECT 3.5950 1.0500 3.9950 1.1500 ;
      RECT 0.3600 1.6250 0.4500 1.9550 ;
      RECT 0.1000 0.4700 0.1900 0.8100 ;
      RECT 0.8800 1.6250 0.9700 1.9550 ;
      RECT 1.4000 1.6250 1.4900 1.9600 ;
      RECT 1.1400 0.4700 1.2300 0.8100 ;
      RECT 0.3600 1.5350 1.8250 1.6250 ;
      RECT 1.7350 1.3500 1.8250 1.5350 ;
      RECT 1.7350 0.9000 1.8250 1.2500 ;
      RECT 0.1000 0.8100 1.8250 0.9000 ;
      RECT 2.5400 1.1500 2.6400 1.2500 ;
      RECT 2.5400 1.0500 2.9500 1.1500 ;
      RECT 3.5950 1.1500 3.6950 1.2500 ;
  END
END AO21B_X6M_A12TH

MACRO AO21_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 0.8700 0.3200 0.9700 0.5600 ;
        RECT 0.0950 0.3200 0.1850 0.7200 ;
        RECT 0.8700 0.5600 1.2800 0.6600 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.3550 1.7500 0.4450 2.0800 ;
        RECT 1.1550 1.5250 1.2450 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.9050 1.5500 1.5000 ;
        RECT 1.4100 1.5000 1.5500 1.9300 ;
        RECT 1.4100 0.4950 1.5500 0.9050 ;
    END
    ANTENNADIFFAREA 0.142625 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.2500 0.3000 1.4000 ;
        RECT 0.0500 1.0800 0.1500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A1

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6800 1.0500 1.1000 1.1500 ;
    END
    ANTENNAGATEAREA 0.0381 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 0.9900 0.5600 1.4000 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A0
  OBS
    LAYER M1 ;
      RECT 0.0950 1.5200 0.7050 1.6100 ;
      RECT 0.6150 1.6100 0.7050 1.9500 ;
      RECT 0.0950 1.6100 0.1850 1.9500 ;
      RECT 0.8900 1.3150 1.3050 1.4050 ;
      RECT 1.2150 0.9000 1.3050 1.3150 ;
      RECT 0.6800 0.8100 1.3050 0.9000 ;
      RECT 0.8900 1.4050 0.9800 1.9400 ;
      RECT 0.6800 0.7200 0.7700 0.8100 ;
      RECT 0.5850 0.5100 0.7700 0.7200 ;
  END
END AO21_X0P5M_A12TH

MACRO ADDF_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.7150 ;
        RECT 0.6200 0.3200 0.7200 0.5600 ;
        RECT 2.1550 0.3200 2.2550 0.6300 ;
        RECT 4.6000 0.3200 4.7000 0.6500 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7250 1.1000 2.1600 1.1500 ;
        RECT 1.4400 1.0600 2.1600 1.1000 ;
        RECT 0.7250 1.1500 1.5400 1.2000 ;
        RECT 1.4400 1.0500 3.7200 1.0600 ;
        RECT 3.6200 1.0600 3.7200 1.1500 ;
        RECT 2.0600 0.9600 3.7200 1.0500 ;
    END
    ANTENNAGATEAREA 0.3402 ;
  END A

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4050 1.4450 3.5900 1.5550 ;
        RECT 3.4050 1.2500 3.5150 1.4450 ;
        RECT 2.2550 1.1900 3.5150 1.2500 ;
        RECT 2.2550 1.2500 2.9000 1.2900 ;
        RECT 2.8000 1.1500 3.5150 1.1900 ;
    END
    ANTENNAGATEAREA 0.2466 ;
  END CI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 3.9700 1.8950 4.1400 2.0800 ;
        RECT 1.1450 1.8000 1.2450 2.0800 ;
        RECT 2.6750 1.8000 2.7750 2.0800 ;
        RECT 2.1550 1.7700 2.2550 2.0800 ;
        RECT 4.6000 1.6050 4.7000 2.0800 ;
        RECT 0.6100 1.5600 0.7100 2.0800 ;
        RECT 0.0900 1.4950 0.1900 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.8700 3.9500 1.2500 ;
        RECT 1.0900 0.8500 3.9500 0.8700 ;
        RECT 1.0900 0.8700 1.9500 0.9500 ;
        RECT 1.8500 0.7700 3.9500 0.8500 ;
        RECT 1.0900 0.9500 1.3000 1.0100 ;
    END
    ANTENNAGATEAREA 0.3402 ;
  END B

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9100 4.5500 1.2900 ;
        RECT 4.3400 1.2900 4.5500 1.3900 ;
        RECT 4.3400 0.8100 4.5500 0.9100 ;
        RECT 4.3400 1.3900 4.4400 1.8300 ;
        RECT 4.3400 0.5300 4.4400 0.8100 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END S

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.2500 ;
        RECT 0.0500 1.2500 0.4500 1.3500 ;
        RECT 0.0500 0.8500 0.4500 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7200 ;
        RECT 0.3500 0.4200 0.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END CO
  OBS
    LAYER M1 ;
      RECT 2.4150 1.5900 3.0650 1.6800 ;
      RECT 2.9650 1.6800 3.0650 1.9900 ;
      RECT 2.4150 1.6800 2.5150 1.9900 ;
      RECT 2.3600 0.4800 3.1300 0.5700 ;
      RECT 0.5400 1.4300 3.1050 1.4700 ;
      RECT 0.5400 1.3800 3.2250 1.4300 ;
      RECT 3.0150 1.3400 3.2250 1.3800 ;
      RECT 0.5400 1.1500 0.6300 1.3800 ;
      RECT 0.3000 1.0500 0.6300 1.1500 ;
      RECT 0.5400 0.7500 0.6300 1.0500 ;
      RECT 1.5700 1.4700 1.7400 1.6850 ;
      RECT 0.5400 0.6600 1.7400 0.7500 ;
      RECT 3.2350 1.6800 4.1900 1.7700 ;
      RECT 4.1000 1.1300 4.1900 1.6800 ;
      RECT 4.1000 1.0300 4.3000 1.1300 ;
      RECT 4.1000 0.6600 4.1900 1.0300 ;
      RECT 3.2250 0.5700 4.1900 0.6600 ;
      RECT 3.2350 1.7700 3.4050 1.9700 ;
      RECT 0.8900 1.5900 1.4650 1.6800 ;
      RECT 1.3750 1.6800 1.4650 1.8300 ;
      RECT 1.3750 1.8300 2.0000 1.9200 ;
      RECT 1.8300 1.6150 2.0000 1.8300 ;
      RECT 0.8900 1.6800 0.9800 1.9800 ;
      RECT 0.8300 0.4800 2.0300 0.5700 ;
  END
END ADDF_X1P4M_A12TH

MACRO ADDF_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0900 0.3200 0.1900 0.6100 ;
        RECT 0.6200 0.3200 0.7200 0.5650 ;
        RECT 2.1550 0.3200 2.2550 0.6300 ;
        RECT 4.6000 0.3200 4.7000 0.6300 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 3.9700 1.8950 4.1400 2.0800 ;
        RECT 0.6100 1.8350 0.7100 2.0800 ;
        RECT 1.1450 1.8000 1.2450 2.0800 ;
        RECT 2.6750 1.8000 2.7750 2.0800 ;
        RECT 0.0900 1.7700 0.1900 2.0800 ;
        RECT 2.1550 1.7700 2.2550 2.0800 ;
        RECT 4.6000 1.7700 4.7000 2.0800 ;
    END
  END VDD

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9500 0.1500 1.2500 ;
        RECT 0.0500 1.2500 0.4500 1.3500 ;
        RECT 0.0500 0.8500 0.4500 0.9500 ;
        RECT 0.3500 1.3500 0.4500 1.7200 ;
        RECT 0.3500 0.4850 0.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END CO

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.9500 4.5500 1.2900 ;
        RECT 4.3400 1.2900 4.5500 1.3900 ;
        RECT 4.3400 0.8500 4.5500 0.9500 ;
        RECT 4.3400 1.3900 4.4400 1.7300 ;
        RECT 4.3400 0.4850 4.4400 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END S

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.8700 3.9500 1.1900 ;
        RECT 1.0900 0.8500 3.9500 0.8700 ;
        RECT 1.0900 0.8700 1.9500 0.9500 ;
        RECT 1.8500 0.7700 3.9500 0.8500 ;
        RECT 1.0900 0.9500 1.3000 1.0100 ;
    END
    ANTENNAGATEAREA 0.3483 ;
  END B

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4050 1.4450 3.5900 1.5550 ;
        RECT 3.4050 1.2500 3.5150 1.4450 ;
        RECT 2.2550 1.1900 3.5150 1.2500 ;
        RECT 2.2550 1.2500 2.9000 1.2900 ;
        RECT 2.8000 1.1500 3.5150 1.1900 ;
    END
    ANTENNAGATEAREA 0.2547 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7250 1.1000 2.1600 1.1500 ;
        RECT 1.4450 1.0600 2.1600 1.1000 ;
        RECT 0.7250 1.1500 1.5450 1.2000 ;
        RECT 1.4450 1.0500 3.7200 1.0600 ;
        RECT 3.6200 1.0600 3.7200 1.1500 ;
        RECT 2.0600 0.9600 3.7200 1.0500 ;
    END
    ANTENNAGATEAREA 0.3483 ;
  END A
  OBS
    LAYER M1 ;
      RECT 2.4150 1.5900 3.0650 1.6800 ;
      RECT 2.9650 1.6800 3.0650 1.9900 ;
      RECT 2.4150 1.6800 2.5150 1.9900 ;
      RECT 2.3600 0.4800 3.1300 0.5700 ;
      RECT 0.5400 1.4300 3.1050 1.4700 ;
      RECT 0.5400 1.3800 3.2250 1.4300 ;
      RECT 3.0150 1.3400 3.2250 1.3800 ;
      RECT 0.5400 1.1500 0.6300 1.3800 ;
      RECT 0.3000 1.0500 0.6300 1.1500 ;
      RECT 0.5400 0.7500 0.6300 1.0500 ;
      RECT 1.5700 1.4700 1.7400 1.6850 ;
      RECT 0.5400 0.6600 1.7400 0.7500 ;
      RECT 3.2350 1.6800 4.1900 1.7700 ;
      RECT 4.1000 1.1500 4.1900 1.6800 ;
      RECT 4.1000 1.0500 4.3000 1.1500 ;
      RECT 4.1000 0.6600 4.1900 1.0500 ;
      RECT 3.2250 0.5700 4.1900 0.6600 ;
      RECT 3.2350 1.7700 3.4050 1.9700 ;
      RECT 0.8900 1.5900 1.4650 1.6800 ;
      RECT 1.3750 1.6800 1.4650 1.8300 ;
      RECT 1.3750 1.8300 2.0000 1.9200 ;
      RECT 1.8300 1.6150 2.0000 1.8300 ;
      RECT 0.8900 1.6800 0.9800 1.9800 ;
      RECT 0.8300 0.4800 2.0300 0.5700 ;
  END
END ADDF_X2M_A12TH

MACRO ADDH_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.6450 0.3200 ;
        RECT 0.3550 0.3200 0.4450 0.7000 ;
        RECT 1.2750 0.3200 1.4450 0.7050 ;
        RECT 2.1000 0.3200 2.1900 0.6500 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5100 1.2500 1.2500 1.3500 ;
        RECT 1.1600 1.1550 1.2500 1.2500 ;
        RECT 0.5100 1.1400 0.6000 1.2500 ;
    END
    ANTENNAGATEAREA 0.1242 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.0650 0.9900 1.1500 ;
        RECT 0.7700 0.9750 1.5100 1.0650 ;
        RECT 1.4200 1.0650 1.5100 1.1450 ;
    END
    ANTENNAGATEAREA 0.1242 ;
  END A

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.4900 0.1700 1.7200 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END CO

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2500 0.9500 2.3500 1.2700 ;
        RECT 2.2500 1.2700 2.4550 1.3700 ;
        RECT 2.2500 0.8500 2.4550 0.9500 ;
        RECT 2.3550 1.3700 2.4550 1.7200 ;
        RECT 2.3550 0.5050 2.4550 0.8500 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.6450 2.7200 ;
        RECT 2.0400 1.7600 2.1300 2.0800 ;
        RECT 0.3400 1.6550 0.4300 2.0800 ;
        RECT 0.9600 1.6400 1.0500 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0550 0.7950 1.6650 0.8850 ;
      RECT 1.5750 0.4100 1.6650 0.7950 ;
      RECT 1.0550 0.4100 1.1450 0.7950 ;
      RECT 0.3300 1.4600 1.4850 1.5500 ;
      RECT 1.3950 1.3800 1.4850 1.4600 ;
      RECT 1.3950 1.2900 1.7400 1.3800 ;
      RECT 1.6500 1.1150 1.7400 1.2900 ;
      RECT 0.3300 1.2100 0.4200 1.4600 ;
      RECT 0.2750 1.0000 0.4200 1.2100 ;
      RECT 0.3150 0.8850 0.4200 1.0000 ;
      RECT 0.6150 1.5500 0.7050 1.8900 ;
      RECT 0.3150 0.7950 0.8950 0.8850 ;
      RECT 0.8050 0.4500 0.8950 0.7950 ;
      RECT 1.8350 1.0750 2.1600 1.1650 ;
      RECT 1.5750 1.5850 1.6650 1.9450 ;
      RECT 1.5750 1.4950 1.9250 1.5850 ;
      RECT 1.8350 1.1650 1.9250 1.4950 ;
      RECT 1.8350 0.4100 1.9250 1.0750 ;
  END
END ADDH_X1M_A12TH

MACRO ADDH_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.8450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.7950 ;
        RECT 0.5400 0.3200 0.7500 0.5400 ;
        RECT 1.1350 0.3200 1.2250 0.4600 ;
        RECT 2.3700 0.3200 2.4600 0.4900 ;
    END
  END VSS

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.4500 0.4300 1.5500 ;
        RECT 0.3400 1.5500 0.4300 1.8700 ;
        RECT 0.0500 0.9850 0.1500 1.4500 ;
        RECT 0.0500 0.8850 0.4300 0.9850 ;
        RECT 0.3400 0.5200 0.4300 0.8850 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END S

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7850 0.8100 0.9900 0.9500 ;
        RECT 0.7850 0.9500 0.8750 1.3950 ;
        RECT 0.7850 1.3950 0.9500 1.4850 ;
        RECT 0.8600 1.4850 0.9500 1.5900 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END CO

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4800 1.0500 2.3950 1.1600 ;
    END
    ANTENNAGATEAREA 0.1608 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2600 1.2500 2.6350 1.3600 ;
        RECT 1.2600 1.1900 1.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.1608 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.8450 2.7200 ;
        RECT 1.1300 1.9900 1.2200 2.0800 ;
        RECT 1.6500 1.9900 1.7400 2.0800 ;
        RECT 0.6000 1.8650 0.6900 2.0800 ;
        RECT 2.6200 1.7900 2.7100 2.0800 ;
        RECT 0.0800 1.6550 0.1700 2.0800 ;
        RECT 1.9000 1.6300 1.9900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0600 1.5000 1.5400 1.5900 ;
      RECT 1.2800 0.8700 2.1550 0.9600 ;
      RECT 1.5950 0.7100 1.6850 0.8700 ;
      RECT 1.0600 1.0100 1.3700 1.1000 ;
      RECT 1.2800 0.9600 1.3700 1.0100 ;
      RECT 1.0600 1.3050 1.1500 1.5000 ;
      RECT 0.9650 1.1000 1.1500 1.3050 ;
      RECT 1.6900 1.4500 2.2500 1.5400 ;
      RECT 2.1600 1.5400 2.2500 1.9400 ;
      RECT 1.3450 0.4800 2.0000 0.5700 ;
      RECT 0.8950 1.7750 1.7800 1.8650 ;
      RECT 1.6900 1.5400 1.7800 1.7750 ;
      RECT 0.6050 0.6300 1.4350 0.7200 ;
      RECT 1.3450 0.5700 1.4350 0.6300 ;
      RECT 0.8950 1.7700 0.9850 1.7750 ;
      RECT 0.6050 1.6800 0.9850 1.7700 ;
      RECT 0.6050 1.3000 0.6950 1.6800 ;
      RECT 0.3000 1.2100 0.6950 1.3000 ;
      RECT 0.6050 0.7200 0.6950 1.2100 ;
      RECT 2.6300 0.7000 2.7200 0.7800 ;
      RECT 2.1100 0.6100 2.7200 0.7000 ;
      RECT 2.6300 0.4100 2.7200 0.6100 ;
      RECT 2.1100 0.4900 2.2000 0.6100 ;
  END
END ADDH_X1P4M_A12TH

MACRO ADDH_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6650 ;
        RECT 0.6000 0.3200 0.6900 0.4800 ;
        RECT 1.2600 0.3200 1.3500 0.6600 ;
        RECT 2.1600 0.3200 2.2500 0.7350 ;
        RECT 2.9700 0.3200 3.0600 0.6000 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8050 0.9500 1.7200 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END CO

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5450 1.2400 2.9050 1.3300 ;
        RECT 1.5450 1.3300 1.9150 1.3500 ;
        RECT 2.8150 1.0500 2.9050 1.2400 ;
    END
    ANTENNAGATEAREA 0.2136 ;
  END A

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.2500 0.4300 1.3500 ;
        RECT 0.3400 1.3500 0.4300 1.7200 ;
        RECT 0.0450 0.9550 0.1350 1.2500 ;
        RECT 0.0450 0.8650 0.4300 0.9550 ;
        RECT 0.3400 0.5200 0.4300 0.8650 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END S

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.5400 2.5500 1.7000 ;
        RECT 2.4500 1.7000 3.2850 1.7200 ;
        RECT 1.2800 1.4400 2.5500 1.5400 ;
        RECT 2.4500 1.7200 3.0100 1.8000 ;
        RECT 2.9100 1.6200 3.2850 1.7000 ;
        RECT 1.2800 1.3450 1.3700 1.4400 ;
        RECT 3.1950 1.0050 3.2850 1.6200 ;
    END
    ANTENNAGATEAREA 0.2136 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 2.1600 1.9400 2.2500 2.0800 ;
        RECT 2.4200 1.9400 2.5100 2.0800 ;
        RECT 1.1200 1.8200 1.2100 2.0800 ;
        RECT 1.6400 1.8200 1.7300 2.0800 ;
        RECT 3.2300 1.8200 3.3200 2.0800 ;
        RECT 0.0800 1.7700 0.1700 2.0800 ;
        RECT 0.6000 1.7700 0.6900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.0400 1.0600 2.6250 1.1500 ;
      RECT 1.0400 1.6400 1.9900 1.7300 ;
      RECT 1.9000 1.7300 1.9900 1.9100 ;
      RECT 1.7100 0.6800 1.8000 1.0600 ;
      RECT 1.0400 1.1500 1.1400 1.6400 ;
      RECT 1.3800 1.7300 1.4700 1.9050 ;
      RECT 2.6700 1.4200 3.1050 1.5100 ;
      RECT 3.0150 0.9600 3.1050 1.4200 ;
      RECT 1.9600 0.8700 3.1050 0.9600 ;
      RECT 1.0600 0.7000 1.1500 0.8550 ;
      RECT 0.6500 0.6100 1.1500 0.7000 ;
      RECT 0.6500 0.7000 0.7400 1.0650 ;
      RECT 0.2450 1.0650 0.7400 1.1550 ;
      RECT 1.9600 0.5700 2.0500 0.8700 ;
      RECT 1.4600 0.4800 2.0500 0.5700 ;
      RECT 1.4600 0.5700 1.5500 0.8550 ;
      RECT 1.0600 0.8550 1.5500 0.9450 ;
      RECT 2.4200 0.4750 2.5100 0.8700 ;
      RECT 2.7100 0.6900 3.3200 0.7800 ;
      RECT 3.2300 0.4100 3.3200 0.6900 ;
      RECT 2.7100 0.4100 2.8000 0.6900 ;
  END
END ADDH_X2M_A12TH

MACRO AND2_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.6950 0.3200 0.7950 0.5600 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5600 1.3950 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0100 0.3500 1.3950 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.6900 1.1500 1.7800 ;
        RECT 0.9800 1.7800 1.1500 1.8800 ;
        RECT 1.0100 0.5900 1.1500 0.6900 ;
        RECT 0.9800 1.8800 1.0800 1.9750 ;
        RECT 1.0100 0.4350 1.1100 0.5900 ;
    END
    ANTENNADIFFAREA 0.167075 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.7200 1.8700 0.8200 2.0800 ;
        RECT 0.1200 1.6800 0.2200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3800 1.5000 0.9500 1.6000 ;
      RECT 0.8500 0.9000 0.9500 1.5000 ;
      RECT 0.1200 0.8000 0.9500 0.9000 ;
      RECT 0.3800 1.6000 0.4800 1.8500 ;
      RECT 0.1200 0.5550 0.2200 0.8000 ;
  END
END AND2_X0P5M_A12TH

MACRO AND2_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.7050 0.3200 0.8050 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.7200 1.7500 0.8200 2.0800 ;
        RECT 0.1200 1.5550 0.2200 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5800 1.3500 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.8750 1.1500 1.5400 ;
        RECT 0.9800 1.5400 1.1500 1.6400 ;
        RECT 0.9800 0.7750 1.1500 0.8750 ;
        RECT 0.9800 1.6400 1.0800 1.9500 ;
        RECT 0.9800 0.4400 1.0800 0.7750 ;
    END
    ANTENNADIFFAREA 0.236775 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.9900 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.3800 1.5300 0.8750 1.6300 ;
      RECT 0.7750 0.8900 0.8750 1.5300 ;
      RECT 0.1200 0.7900 0.8750 0.8900 ;
      RECT 0.3800 1.6300 0.4800 1.7450 ;
      RECT 0.1200 0.5950 0.2200 0.7900 ;
  END
END AND2_X0P7M_A12TH

MACRO AND2_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.1200 0.3200 0.2200 0.6350 ;
        RECT 1.0600 0.3200 1.1600 0.5900 ;
        RECT 2.0000 0.3200 2.1000 0.5900 ;
        RECT 2.9850 0.3200 3.0850 0.5900 ;
        RECT 3.5500 0.3200 3.6500 0.6350 ;
        RECT 4.0700 0.3200 4.1700 0.6350 ;
        RECT 4.5900 0.3200 4.6900 0.6350 ;
        RECT 5.1100 0.3200 5.2100 0.6350 ;
        RECT 5.6300 0.3200 5.7300 0.6350 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8200 0.9300 5.9950 1.2800 ;
        RECT 3.2600 1.2800 5.9950 1.4400 ;
        RECT 3.2600 0.7700 5.9950 0.9300 ;
        RECT 3.2600 1.4400 3.4200 1.7400 ;
        RECT 3.7800 1.4400 3.9400 1.7450 ;
        RECT 4.3000 1.4400 4.4600 1.7450 ;
        RECT 4.8200 1.4400 4.9800 1.7450 ;
        RECT 5.3400 1.4400 5.5000 1.7450 ;
        RECT 5.8600 1.4400 5.9950 1.7450 ;
        RECT 3.2600 0.4700 3.4200 0.7700 ;
        RECT 3.7800 0.4700 3.9400 0.7700 ;
        RECT 4.3000 0.4700 4.4600 0.7700 ;
        RECT 4.8200 0.4700 4.9800 0.7700 ;
        RECT 5.3400 0.4700 5.5000 0.7700 ;
        RECT 5.8600 0.4700 5.9950 0.7700 ;
    END
    ANTENNADIFFAREA 1.958125 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.2900 2.9500 1.3900 ;
        RECT 1.0300 1.3900 2.1850 1.4250 ;
        RECT 0.2400 1.0400 0.3400 1.2900 ;
        RECT 2.8400 1.0200 2.9500 1.2900 ;
    END
    ANTENNAGATEAREA 0.4284 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4600 1.0500 2.7200 1.1500 ;
    END
    ANTENNAGATEAREA 0.4284 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.3900 1.7700 0.4900 2.0800 ;
        RECT 0.9100 1.7700 1.0100 2.0800 ;
        RECT 1.4300 1.7700 1.5300 2.0800 ;
        RECT 1.9500 1.7700 2.0500 2.0800 ;
        RECT 2.4700 1.7700 2.5700 2.0800 ;
        RECT 3.0150 1.7700 3.1150 2.0800 ;
        RECT 3.5500 1.7700 3.6500 2.0800 ;
        RECT 4.0700 1.7700 4.1700 2.0800 ;
        RECT 4.5900 1.7700 4.6900 2.0800 ;
        RECT 5.1100 1.7700 5.2100 2.0800 ;
        RECT 5.6300 1.7700 5.7300 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 3.0400 1.0550 4.8300 1.1550 ;
      RECT 0.6500 1.6450 0.7500 1.9550 ;
      RECT 0.5900 0.4200 0.6900 0.7100 ;
      RECT 1.1700 1.6450 1.2700 1.9550 ;
      RECT 1.6900 1.6450 1.7900 1.9550 ;
      RECT 1.5300 0.4200 1.6300 0.7100 ;
      RECT 2.2100 1.6450 2.3100 1.9550 ;
      RECT 2.7300 1.6450 2.8300 1.9550 ;
      RECT 2.4700 0.4200 2.5700 0.7100 ;
      RECT 0.6500 1.5450 3.1400 1.6450 ;
      RECT 3.0400 1.1550 3.1400 1.5450 ;
      RECT 3.0400 0.8100 3.1400 1.0550 ;
      RECT 0.5900 0.7100 3.1400 0.8100 ;
  END
END AND2_X11M_A12TH

MACRO AND2_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.2450 0.3200 ;
        RECT 0.7050 0.3200 0.8050 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0000 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0500 0.9100 1.1500 1.2900 ;
        RECT 0.9800 1.2900 1.1500 1.3900 ;
        RECT 0.9800 0.8100 1.1500 0.9100 ;
        RECT 0.9800 1.3900 1.0800 1.7200 ;
        RECT 0.9800 0.4800 1.0800 0.8100 ;
    END
    ANTENNADIFFAREA 0.333125 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5800 1.3500 ;
    END
    ANTENNAGATEAREA 0.0414 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.2450 2.7200 ;
        RECT 0.7200 1.7700 0.8200 2.0800 ;
        RECT 0.1200 1.5800 0.2200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3250 1.5650 0.8600 1.6650 ;
      RECT 0.7600 0.8800 0.8600 1.5650 ;
      RECT 0.1200 0.7800 0.8600 0.8800 ;
      RECT 0.1200 0.4900 0.2200 0.7800 ;
  END
END AND2_X1M_A12TH

MACRO AND2_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6300 0.3200 0.7300 0.6450 ;
        RECT 1.1900 0.3200 1.2900 0.8000 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1900 1.7200 1.2900 2.0800 ;
        RECT 0.6550 1.7100 0.7550 2.0800 ;
        RECT 0.1200 1.4900 0.2200 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.5800 1.3500 ;
    END
    ANTENNAGATEAREA 0.0567 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0200 1.3500 1.4500 ;
        RECT 0.9300 1.4500 1.3500 1.5500 ;
        RECT 0.9300 0.9200 1.3500 1.0200 ;
        RECT 0.9300 1.5500 1.0300 1.9350 ;
        RECT 0.9300 0.5000 1.0300 0.9200 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0567 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.7000 1.1800 1.1600 1.2700 ;
      RECT 0.3800 1.5000 0.8000 1.6000 ;
      RECT 0.7000 1.2700 0.8000 1.5000 ;
      RECT 0.7000 0.8850 0.8000 1.1800 ;
      RECT 0.1200 0.7850 0.8000 0.8850 ;
      RECT 0.3800 1.6000 0.4800 1.9350 ;
      RECT 0.1200 0.4550 0.2200 0.7850 ;
  END
END AND2_X1P4M_A12TH

MACRO AND2_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.6300 0.3200 0.7300 0.6400 ;
        RECT 1.1900 0.3200 1.2900 0.6350 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 1.0100 0.5800 1.3900 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 1.1900 1.7700 1.2900 2.0800 ;
        RECT 0.6550 1.6700 0.7550 2.0800 ;
        RECT 0.1200 1.4800 0.2200 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9500 1.3500 1.4500 ;
        RECT 0.9300 1.4500 1.3500 1.5500 ;
        RECT 0.9300 0.8500 1.3500 0.9500 ;
        RECT 0.9300 1.5500 1.0300 1.8900 ;
        RECT 0.9300 0.4700 1.0300 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0050 0.3500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0762 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.7100 1.0600 1.1600 1.1500 ;
      RECT 0.3800 1.4800 0.8100 1.5800 ;
      RECT 0.7100 1.1500 0.8100 1.4800 ;
      RECT 0.7100 0.8850 0.8100 1.0600 ;
      RECT 0.1200 0.7850 0.8100 0.8850 ;
      RECT 0.3800 1.5800 0.4800 1.8800 ;
      RECT 0.1200 0.4550 0.2200 0.7850 ;
  END
END AND2_X2M_A12TH

MACRO AND2_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.0450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6550 ;
        RECT 0.8550 0.3200 0.9550 0.6550 ;
        RECT 1.8250 0.3200 1.9250 0.8250 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9900 1.2500 1.7500 1.3500 ;
        RECT 1.6500 1.3500 1.7500 1.5200 ;
        RECT 0.9900 1.0100 1.0900 1.2500 ;
    END
    ANTENNAGATEAREA 0.117 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2350 1.0500 1.7050 1.1500 ;
    END
    ANTENNAGATEAREA 0.117 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0700 1.2500 0.6950 1.3500 ;
        RECT 0.0700 1.3500 0.1700 1.7200 ;
        RECT 0.5950 1.3500 0.6950 1.7200 ;
        RECT 0.0700 0.9400 0.1700 1.2500 ;
        RECT 0.0700 0.8400 0.6950 0.9400 ;
        RECT 0.0700 0.5100 0.1700 0.8400 ;
        RECT 0.5950 0.5100 0.6950 0.8400 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.0450 2.7200 ;
        RECT 0.3350 1.7700 0.4350 2.0800 ;
        RECT 0.8550 1.7200 0.9550 2.0800 ;
        RECT 1.4000 1.7200 1.5000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.8100 0.8000 1.4750 0.8900 ;
      RECT 1.3750 0.4700 1.4750 0.8000 ;
      RECT 1.1450 1.5700 1.2350 1.9000 ;
      RECT 0.8100 1.4800 1.2350 1.5700 ;
      RECT 0.8100 1.1500 0.9000 1.4800 ;
      RECT 0.2950 1.0600 0.9000 1.1500 ;
      RECT 0.8100 0.8900 0.9000 1.0600 ;
  END
END AND2_X3M_A12TH

MACRO AND2_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.4450 0.3200 ;
        RECT 0.1500 0.3200 0.2500 0.6400 ;
        RECT 1.1300 0.3200 1.2300 0.6400 ;
        RECT 1.6900 0.3200 1.7900 0.6350 ;
        RECT 2.2100 0.3200 2.3100 0.6350 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 1.0500 1.0850 1.1500 ;
        RECT 0.9850 1.1500 1.0850 1.3600 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.4450 2.7200 ;
        RECT 0.6200 1.7900 0.7200 2.0800 ;
        RECT 1.1550 1.7900 1.2550 2.0800 ;
        RECT 0.1000 1.7700 0.2000 2.0800 ;
        RECT 1.6900 1.7700 1.7900 2.0800 ;
        RECT 2.2100 1.7700 2.3100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9100 2.1500 1.4500 ;
        RECT 1.4300 1.4500 2.1500 1.5500 ;
        RECT 1.4300 0.8100 2.1500 0.9100 ;
        RECT 1.4300 1.5500 1.5300 1.8600 ;
        RECT 1.9500 1.5500 2.0500 1.8600 ;
        RECT 1.4300 0.4700 1.5300 0.8100 ;
        RECT 1.9500 0.4700 2.0500 0.8100 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4800 1.2450 0.8750 1.3550 ;
    END
    ANTENNAGATEAREA 0.1524 ;
  END A
  OBS
    LAYER M1 ;
      RECT 1.2050 1.0550 1.9300 1.1550 ;
      RECT 0.3600 1.7000 0.4600 1.9850 ;
      RECT 0.8800 1.7000 0.9800 1.9850 ;
      RECT 0.6200 0.4400 0.7200 0.8400 ;
      RECT 0.3600 1.6000 1.3050 1.7000 ;
      RECT 1.2050 1.1550 1.3050 1.6000 ;
      RECT 1.2050 0.9400 1.3050 1.0550 ;
      RECT 0.6200 0.8400 1.3050 0.9400 ;
  END
END AND2_X4M_A12TH

MACRO AND2_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.5900 0.3200 0.6900 0.5600 ;
        RECT 1.5750 0.3200 1.6750 0.5600 ;
        RECT 2.1400 0.3200 2.2400 0.6350 ;
        RECT 2.6600 0.3200 2.7600 0.6350 ;
        RECT 3.1800 0.3200 3.2800 0.6350 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9200 1.0500 1.2900 1.1500 ;
        RECT 0.9200 1.1500 1.0200 1.2850 ;
        RECT 0.2400 1.2850 1.0200 1.3850 ;
        RECT 0.2400 1.0450 0.3500 1.2850 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0500 0.9050 3.1500 1.2900 ;
        RECT 1.8800 1.2900 3.1500 1.3900 ;
        RECT 1.8800 0.8050 3.1500 0.9050 ;
        RECT 1.8800 1.3900 1.9800 1.7400 ;
        RECT 2.4000 1.3900 2.5000 1.7450 ;
        RECT 2.9200 1.3900 3.0200 1.7450 ;
        RECT 1.8800 0.4700 1.9800 0.8050 ;
        RECT 2.4000 0.4700 2.5000 0.8050 ;
        RECT 2.9200 0.4700 3.0200 0.8050 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4550 1.0500 0.8250 1.1500 ;
        RECT 0.7250 0.9500 0.8250 1.0500 ;
        RECT 0.7250 0.8500 1.5500 0.9500 ;
        RECT 1.4500 0.9500 1.5500 1.3050 ;
    END
    ANTENNAGATEAREA 0.2316 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.5400 1.7700 0.6400 2.0800 ;
        RECT 1.0600 1.7700 1.1600 2.0800 ;
        RECT 1.6050 1.7700 1.7050 2.0800 ;
        RECT 2.1400 1.7700 2.2400 2.0800 ;
        RECT 2.6600 1.7700 2.7600 2.0800 ;
        RECT 3.1800 1.7700 3.2800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.6500 1.0550 2.7100 1.1550 ;
      RECT 0.8000 1.5450 1.7500 1.6450 ;
      RECT 1.6500 1.1550 1.7500 1.5450 ;
      RECT 1.6500 0.7500 1.7500 1.0550 ;
      RECT 0.0850 0.6500 1.7500 0.7500 ;
      RECT 0.0850 0.4100 0.2550 0.6500 ;
      RECT 1.3200 1.6450 1.4200 1.9550 ;
      RECT 1.0250 0.4100 1.1950 0.6500 ;
      RECT 0.8000 1.6450 0.9000 1.9550 ;
  END
END AND2_X6M_A12TH

MACRO AND2_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6500 ;
        RECT 0.9800 0.3200 1.0700 0.6500 ;
        RECT 1.9350 0.3200 2.0250 0.6500 ;
        RECT 2.4700 0.3200 2.5600 0.6500 ;
        RECT 2.9900 0.3200 3.0800 0.6500 ;
        RECT 3.5100 0.3200 3.6000 0.6500 ;
        RECT 4.0300 0.3200 4.1200 0.6500 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4350 1.0500 1.6950 1.1250 ;
        RECT 0.6100 1.1250 1.6950 1.1500 ;
        RECT 0.4350 1.0250 0.7650 1.0500 ;
    END
    ANTENNAGATEAREA 0.3087 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2550 1.2500 1.8950 1.3500 ;
        RECT 0.2550 1.3500 1.1800 1.3550 ;
        RECT 0.2550 1.2150 0.3450 1.2500 ;
        RECT 1.8050 1.1350 1.8950 1.2500 ;
        RECT 0.2550 1.3550 0.3450 1.4150 ;
    END
    ANTENNAGATEAREA 0.3087 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 1.9500 1.7700 2.0400 2.0800 ;
        RECT 2.4700 1.7700 2.5600 2.0800 ;
        RECT 2.9900 1.7700 3.0800 2.0800 ;
        RECT 3.5100 1.7700 3.6000 2.0800 ;
        RECT 4.0300 1.7700 4.1200 2.0800 ;
        RECT 0.3800 1.7500 0.4700 2.0800 ;
        RECT 0.9000 1.7500 0.9900 2.0800 ;
        RECT 1.4200 1.7500 1.5100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8350 0.9650 3.9650 1.4350 ;
        RECT 2.1950 1.4350 3.9650 1.5650 ;
        RECT 2.1900 0.8350 3.9650 0.9650 ;
        RECT 2.1950 1.5650 2.3250 1.8850 ;
        RECT 2.7300 1.5650 2.8200 1.8850 ;
        RECT 3.2500 1.5650 3.3400 1.8850 ;
        RECT 3.7700 1.5650 3.8600 1.8800 ;
        RECT 2.1900 0.4850 2.3200 0.8350 ;
        RECT 2.7300 0.4850 2.8200 0.8350 ;
        RECT 3.2500 0.4850 3.3400 0.8350 ;
        RECT 3.7700 0.4850 3.8600 0.8350 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.9850 1.0900 3.6750 1.1800 ;
      RECT 0.6400 1.5550 0.7300 1.8950 ;
      RECT 0.5300 0.4850 0.6200 0.8250 ;
      RECT 1.1600 1.5550 1.2500 1.8950 ;
      RECT 1.6800 1.5550 1.7700 1.8950 ;
      RECT 1.4700 0.4850 1.5600 0.8250 ;
      RECT 0.6400 1.4650 2.0750 1.5550 ;
      RECT 1.9850 1.1800 2.0750 1.4650 ;
      RECT 1.9850 0.9150 2.0750 1.0900 ;
      RECT 0.5300 0.8250 2.0750 0.9150 ;
  END
END AND2_X8M_A12TH

MACRO AND3_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.8750 0.3200 0.9650 0.9100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 0.9900 0.3500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.6950 0.7550 1.0200 ;
        RECT 0.6500 1.0200 0.8800 1.1100 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 0.7050 1.4050 ;
        RECT 0.4500 1.0800 0.5500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9800 1.3500 1.4100 ;
        RECT 1.1750 1.4100 1.3500 1.5100 ;
        RECT 1.1800 0.8800 1.3500 0.9800 ;
        RECT 1.1750 1.5100 1.2750 1.8400 ;
        RECT 1.1800 0.5100 1.2800 0.8800 ;
    END
    ANTENNADIFFAREA 0.167075 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3800 1.7200 0.4800 2.0800 ;
        RECT 0.9000 1.7200 1.0000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0550 1.5300 1.0700 1.6300 ;
      RECT 0.9700 1.2050 1.0700 1.5300 ;
      RECT 0.9700 1.1150 1.1500 1.2050 ;
      RECT 0.0550 0.7900 0.2750 0.8800 ;
      RECT 0.1850 0.5000 0.2750 0.7900 ;
      RECT 0.1200 1.6300 0.2200 1.8600 ;
      RECT 0.0550 0.8800 0.1450 1.5300 ;
      RECT 0.6400 1.6300 0.7400 1.8600 ;
  END
END AND3_X0P5M_A12TH

MACRO AND3_X0P7M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.8850 0.3200 0.9850 0.9000 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9550 1.3500 1.3450 ;
        RECT 1.1750 1.3450 1.3500 1.4450 ;
        RECT 1.1750 0.8100 1.3500 0.9550 ;
        RECT 1.1750 1.4450 1.2750 1.7750 ;
        RECT 1.1750 0.5100 1.2750 0.8100 ;
    END
    ANTENNADIFFAREA 0.236775 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 0.7050 1.3900 ;
        RECT 0.4500 1.0800 0.5500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.6950 0.7500 1.0700 ;
        RECT 0.6500 1.0700 0.8800 1.1600 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3550 1.4100 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3800 1.7800 0.4800 2.0800 ;
        RECT 0.9000 1.7800 1.0000 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.5450 1.0700 1.6450 ;
      RECT 0.9700 1.2050 1.0700 1.5450 ;
      RECT 0.9700 1.1150 1.1500 1.2050 ;
      RECT 0.0500 0.7900 0.2800 0.8900 ;
      RECT 0.1800 0.4600 0.2800 0.7900 ;
      RECT 0.1200 1.6450 0.2200 1.9300 ;
      RECT 0.0500 0.8900 0.1500 1.5450 ;
      RECT 0.6400 1.6450 0.7400 1.9300 ;
  END
END AND3_X0P7M_A12TH

MACRO AND3_X11M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 9.0450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6300 ;
        RECT 1.3650 0.3200 1.5350 0.5200 ;
        RECT 2.6850 0.3200 2.8550 0.5200 ;
        RECT 4.2450 0.3200 4.4150 0.5200 ;
        RECT 5.8650 0.3200 6.0350 0.5200 ;
        RECT 6.4900 0.3200 6.5800 0.6850 ;
        RECT 7.0100 0.3200 7.1000 0.6850 ;
        RECT 7.5300 0.3200 7.6200 0.6850 ;
        RECT 8.0500 0.3200 8.1400 0.6850 ;
        RECT 8.5700 0.3200 8.6600 0.6850 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3950 1.2600 1.8850 1.3500 ;
        RECT 0.3950 1.3500 0.4850 1.4700 ;
        RECT 0.3950 1.2500 1.7500 1.2600 ;
        RECT 1.6500 0.9900 1.7500 1.2500 ;
        RECT 1.6500 0.9000 3.1800 0.9900 ;
        RECT 2.3400 0.9900 2.4300 1.2600 ;
        RECT 3.0900 0.9900 3.1800 1.2100 ;
        RECT 3.0900 0.8800 3.1800 0.9000 ;
        RECT 2.2200 1.2600 2.4300 1.3500 ;
        RECT 3.0900 0.8700 5.6600 0.8800 ;
        RECT 3.9200 0.8800 4.7800 0.9600 ;
        RECT 5.5700 0.8800 5.6600 1.2100 ;
        RECT 3.0900 0.7900 4.0100 0.8700 ;
        RECT 4.6900 0.7900 5.6600 0.8700 ;
        RECT 3.9200 0.9600 4.0100 1.2100 ;
        RECT 4.5900 0.9600 4.7800 1.1300 ;
    END
    ANTENNAGATEAREA 0.582 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.2500 3.5500 1.5000 ;
        RECT 0.6150 1.5000 5.0350 1.5900 ;
        RECT 3.4500 1.1500 3.6300 1.2500 ;
        RECT 4.9450 1.4900 5.0350 1.5000 ;
        RECT 4.9450 1.4000 5.1400 1.4900 ;
        RECT 5.0500 1.2400 5.1400 1.4000 ;
        RECT 5.0500 1.1500 5.2600 1.2400 ;
    END
    ANTENNAGATEAREA 0.582 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1200 1.2200 4.9600 1.3100 ;
        RECT 4.1200 1.3100 4.4100 1.3200 ;
        RECT 4.1200 1.0900 4.5000 1.2200 ;
        RECT 4.8700 1.0600 4.9600 1.2200 ;
        RECT 3.7400 1.3200 4.4100 1.3500 ;
        RECT 4.8700 0.9700 5.4600 1.0600 ;
        RECT 3.7400 1.3500 4.2450 1.4100 ;
        RECT 3.7400 1.0600 3.8300 1.3200 ;
        RECT 5.3700 1.0600 5.4600 1.3000 ;
        RECT 3.2700 0.9700 3.8300 1.0600 ;
        RECT 5.3700 1.3000 5.8900 1.3900 ;
        RECT 3.2700 1.0600 3.3600 1.3200 ;
        RECT 5.8000 1.0500 5.8900 1.3000 ;
        RECT 2.9100 1.3200 3.3600 1.4100 ;
        RECT 2.9100 1.2000 3.0000 1.3200 ;
        RECT 2.5900 1.1100 3.0000 1.2000 ;
    END
    ANTENNAGATEAREA 0.582 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.1950 1.4200 8.9550 1.5800 ;
        RECT 6.1950 1.5800 6.3550 1.8500 ;
        RECT 6.7150 1.5800 6.8750 1.8500 ;
        RECT 7.2350 1.5800 7.3950 1.8500 ;
        RECT 7.7550 1.5800 7.9150 1.8500 ;
        RECT 8.2750 1.5800 8.4350 1.8500 ;
        RECT 8.7950 1.5800 8.9550 1.8500 ;
        RECT 8.6200 0.9800 8.7800 1.4200 ;
        RECT 6.1950 0.8200 8.9550 0.9800 ;
        RECT 6.1950 0.5400 6.3550 0.8200 ;
        RECT 6.7150 0.5400 6.8750 0.8200 ;
        RECT 7.2350 0.5400 7.3950 0.8200 ;
        RECT 7.7550 0.5400 7.9150 0.8200 ;
        RECT 8.2750 0.5400 8.4350 0.8200 ;
        RECT 8.7950 0.5350 8.9550 0.8200 ;
    END
    ANTENNADIFFAREA 1.885 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 9.0450 2.7200 ;
        RECT 3.2050 1.8750 3.3750 2.0800 ;
        RECT 3.7250 1.8750 3.8950 2.0800 ;
        RECT 4.2450 1.8750 4.4150 2.0800 ;
        RECT 4.7850 1.8750 4.9550 2.0800 ;
        RECT 5.3450 1.8750 5.5150 2.0800 ;
        RECT 5.9250 1.8750 6.0950 2.0800 ;
        RECT 2.7250 1.8000 2.8150 2.0800 ;
        RECT 6.4900 1.7700 6.5800 2.0800 ;
        RECT 7.0100 1.7700 7.1000 2.0800 ;
        RECT 7.5300 1.7700 7.6200 2.0800 ;
        RECT 8.0500 1.7700 8.1400 2.0800 ;
        RECT 8.5700 1.7700 8.6600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 5.9800 1.0800 8.3300 1.1700 ;
      RECT 0.7450 0.4200 0.8350 0.6350 ;
      RECT 0.7450 0.7250 0.8350 0.8500 ;
      RECT 0.7450 0.7000 2.1550 0.7250 ;
      RECT 2.0650 0.7250 2.1550 0.8100 ;
      RECT 2.0650 0.4400 2.1550 0.6100 ;
      RECT 2.9450 1.7700 3.1150 1.9700 ;
      RECT 3.4650 1.7700 3.6350 1.9700 ;
      RECT 3.4650 0.4100 3.6350 0.6100 ;
      RECT 3.9850 1.7700 4.1550 1.9700 ;
      RECT 4.5050 1.7700 4.6750 1.9700 ;
      RECT 5.1250 1.7700 5.2150 1.9850 ;
      RECT 5.1250 1.6150 5.2150 1.6800 ;
      RECT 5.0850 0.4100 5.2550 0.6100 ;
      RECT 5.6450 1.7700 5.7350 1.9850 ;
      RECT 5.6450 1.6150 5.7350 1.6800 ;
      RECT 2.9450 1.6800 6.0700 1.7700 ;
      RECT 5.9800 1.1700 6.0700 1.6800 ;
      RECT 5.9800 0.7000 6.0700 1.0800 ;
      RECT 0.7450 0.6350 6.0700 0.7000 ;
      RECT 2.0650 0.6100 6.0700 0.6350 ;
  END
END AND3_X11M_A12TH

MACRO AND3_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.4450 0.3200 ;
        RECT 0.8850 0.3200 0.9850 0.7450 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3550 1.4100 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6500 0.6950 0.7650 1.0700 ;
        RECT 0.6500 1.0700 0.8800 1.1600 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.2500 0.7050 1.3900 ;
        RECT 0.4500 1.0800 0.5500 1.2500 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 0.9100 1.3500 1.2900 ;
        RECT 1.1750 1.2900 1.3500 1.3900 ;
        RECT 1.1750 0.8100 1.3500 0.9100 ;
        RECT 1.1750 1.3900 1.2750 1.7200 ;
        RECT 1.1750 0.4800 1.2750 0.8100 ;
    END
    ANTENNADIFFAREA 0.333125 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.4450 2.7200 ;
        RECT 0.3450 1.7250 0.5150 2.0800 ;
        RECT 0.8650 1.7250 1.0350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0500 1.5250 1.0700 1.6250 ;
      RECT 0.9700 1.1500 1.0700 1.5250 ;
      RECT 0.9700 1.0600 1.1500 1.1500 ;
      RECT 0.0500 0.7900 0.2800 0.8900 ;
      RECT 0.1800 0.4600 0.2800 0.7900 ;
      RECT 0.1200 1.6300 0.2200 1.8950 ;
      RECT 0.0500 1.6250 0.2200 1.6300 ;
      RECT 0.0500 0.8900 0.1500 1.5250 ;
      RECT 0.6400 1.6250 0.7400 1.8900 ;
  END
END AND3_X1M_A12TH

MACRO AND3_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.8450 0.3200 ;
        RECT 1.0600 0.3200 1.1600 0.7150 ;
        RECT 1.6150 0.3200 1.7050 0.7150 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.9500 1.7500 1.4500 ;
        RECT 1.3500 1.4500 1.7500 1.5500 ;
        RECT 1.3500 0.8500 1.7500 0.9500 ;
        RECT 1.3500 1.5500 1.4500 1.8800 ;
        RECT 1.3500 0.4150 1.4500 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6400 1.0900 0.7550 1.4900 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 0.8800 0.9500 1.1600 ;
        RECT 0.8500 1.1600 1.0150 1.3700 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.0100 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0828 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.8450 2.7200 ;
        RECT 0.5550 1.8600 0.6550 2.0800 ;
        RECT 1.0750 1.8600 1.1750 2.0800 ;
        RECT 1.6200 1.6800 1.7200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1450 1.0700 1.5450 1.2400 ;
      RECT 0.0500 1.5900 1.2450 1.6900 ;
      RECT 1.1450 1.2400 1.2450 1.5900 ;
      RECT 0.2950 1.6900 0.3950 1.9850 ;
      RECT 0.0500 0.7900 0.4550 0.8900 ;
      RECT 0.3550 0.4600 0.4550 0.7900 ;
      RECT 0.0500 0.8900 0.1500 1.5900 ;
      RECT 0.8150 1.6900 0.9150 1.9850 ;
  END
END AND3_X1P4M_A12TH

MACRO AND3_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 2.2450 0.3200 ;
        RECT 0.1150 0.3200 0.2150 0.7750 ;
        RECT 1.4450 0.3200 1.5450 0.6900 ;
        RECT 2.0100 0.3200 2.1100 0.6350 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4350 1.2500 1.1600 1.3500 ;
    END
    ANTENNAGATEAREA 0.1086 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.4500 1.4000 1.5500 ;
        RECT 0.2800 1.5500 0.3950 1.6200 ;
        RECT 1.3000 1.0400 1.4000 1.4500 ;
    END
    ANTENNAGATEAREA 0.1086 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6950 1.0300 1.1100 1.1500 ;
    END
    ANTENNAGATEAREA 0.1086 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 2.2450 2.7200 ;
        RECT 0.8750 1.8400 0.9750 2.0800 ;
        RECT 1.4450 1.8400 1.5450 2.0800 ;
        RECT 2.0100 1.7700 2.1100 2.0800 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0500 0.9500 2.1500 1.2600 ;
        RECT 1.7500 1.2600 2.1500 1.3600 ;
        RECT 1.7500 0.8500 2.1500 0.9500 ;
        RECT 1.7500 1.3600 1.8500 1.7200 ;
        RECT 1.7500 0.4900 1.8500 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 1.5450 1.0600 1.9600 1.1500 ;
      RECT 0.5800 1.6400 1.6450 1.7400 ;
      RECT 1.5450 1.1500 1.6450 1.6400 ;
      RECT 1.5450 0.9100 1.6450 1.0600 ;
      RECT 0.7550 0.8100 1.6450 0.9100 ;
      RECT 0.5800 1.7400 0.7500 1.9900 ;
      RECT 0.7550 0.4600 0.8550 0.8100 ;
      RECT 1.1000 1.7400 1.2700 1.9900 ;
  END
END AND3_X2M_A12TH

MACRO AND3_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.0450 0.3200 ;
        RECT 0.7200 0.3200 0.8100 0.5800 ;
        RECT 2.0500 0.3200 2.1400 0.6500 ;
        RECT 2.5700 0.3200 2.6600 0.6500 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5550 0.8700 2.0200 0.9600 ;
        RECT 0.5550 0.9600 0.9450 1.0200 ;
        RECT 1.9300 0.9600 2.0200 1.1550 ;
        RECT 0.5550 0.8500 0.8550 0.8700 ;
    END
    ANTENNAGATEAREA 0.1608 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0650 1.0900 1.8200 1.1100 ;
        RECT 0.2850 1.1100 1.8200 1.2000 ;
        RECT 1.0650 1.0800 1.5900 1.0900 ;
        RECT 0.7550 1.2000 0.9650 1.2800 ;
        RECT 1.2750 1.0500 1.5900 1.0800 ;
    END
    ANTENNAGATEAREA 0.1608 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.4500 1.2300 1.5500 ;
        RECT 1.1400 1.4200 1.2300 1.4500 ;
        RECT 0.2800 1.3400 0.3700 1.4500 ;
        RECT 1.1400 1.3200 1.5300 1.4200 ;
    END
    ANTENNAGATEAREA 0.1608 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3100 1.4500 2.9200 1.5500 ;
        RECT 2.3100 1.5500 2.4000 1.8800 ;
        RECT 2.8300 1.5500 2.9200 1.8600 ;
        RECT 2.8300 0.9450 2.9200 1.4500 ;
        RECT 2.3100 0.8550 2.9200 0.9450 ;
        RECT 2.3100 0.5050 2.4000 0.8550 ;
        RECT 2.8300 0.5050 2.9200 0.8550 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.0450 2.7200 ;
        RECT 0.4750 1.8250 0.5650 2.0800 ;
        RECT 0.9950 1.8250 1.0850 2.0800 ;
        RECT 1.5150 1.8250 1.6050 2.0800 ;
        RECT 2.0500 1.8250 2.1400 2.0800 ;
        RECT 2.5700 1.7700 2.6600 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.1300 1.0900 2.6050 1.1800 ;
      RECT 0.0800 0.7600 0.1700 1.6400 ;
      RECT 0.0800 0.4100 0.1700 0.6700 ;
      RECT 0.6950 1.7350 0.8650 1.9900 ;
      RECT 1.2150 1.7350 1.3850 1.9900 ;
      RECT 0.0800 0.6700 1.4500 0.7600 ;
      RECT 1.3600 0.7600 1.4500 0.7800 ;
      RECT 1.3600 0.4100 1.4500 0.6700 ;
      RECT 0.0800 1.7300 1.9050 1.7350 ;
      RECT 1.7350 1.7350 1.9050 1.9900 ;
      RECT 0.0800 1.6400 2.2200 1.7300 ;
      RECT 2.1300 1.1800 2.2200 1.6400 ;
  END
END AND3_X3M_A12TH

MACRO AND3_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 3.4450 0.3200 ;
        RECT 0.7450 0.3200 0.8350 0.5800 ;
        RECT 2.1750 0.3200 2.2650 0.6700 ;
        RECT 2.7100 0.3200 2.8000 0.6700 ;
        RECT 3.2300 0.3200 3.3200 0.6700 ;
    END
  END VSS

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4100 0.8500 0.5900 1.0150 ;
        RECT 0.4100 1.0150 0.9000 1.1150 ;
        RECT 0.8100 0.9600 0.9000 1.0150 ;
        RECT 0.8100 0.8700 2.1650 0.9600 ;
        RECT 2.0750 0.9600 2.1650 1.2450 ;
    END
    ANTENNAGATEAREA 0.2079 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3350 1.2500 1.1150 1.3500 ;
        RECT 0.9450 1.3500 1.1150 1.3850 ;
        RECT 1.0150 1.1500 1.1150 1.2500 ;
        RECT 1.0150 1.0500 1.9450 1.1500 ;
        RECT 1.8450 1.1500 1.9450 1.4600 ;
    END
    ANTENNAGATEAREA 0.2079 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2800 1.4850 1.3900 1.5650 ;
        RECT 0.2800 1.5650 0.4900 1.5750 ;
        RECT 0.4000 1.4750 1.6550 1.4850 ;
        RECT 1.2100 1.3850 1.6550 1.4750 ;
    END
    ANTENNAGATEAREA 0.2079 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4500 1.4500 3.1650 1.5500 ;
        RECT 2.4500 1.5500 2.5400 1.8800 ;
        RECT 2.9700 1.5500 3.0600 1.8800 ;
        RECT 3.0750 0.9800 3.1650 1.4500 ;
        RECT 2.4500 0.8900 3.1650 0.9800 ;
        RECT 2.4500 0.5250 2.5400 0.8900 ;
        RECT 2.9700 0.5250 3.0600 0.8900 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 3.4450 2.7200 ;
        RECT 0.5800 1.8600 0.7500 2.0800 ;
        RECT 1.1000 1.8600 1.2700 2.0800 ;
        RECT 1.6200 1.8600 1.7900 2.0800 ;
        RECT 2.1500 1.8600 2.3200 2.0800 ;
        RECT 2.7100 1.7700 2.8000 2.0800 ;
        RECT 3.2300 1.7700 3.3200 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 2.2550 1.0900 2.9850 1.1800 ;
      RECT 0.0800 0.7600 0.1700 1.6650 ;
      RECT 0.0800 0.4100 0.1700 0.6700 ;
      RECT 0.8400 1.7550 1.0100 1.9550 ;
      RECT 1.3600 1.7550 1.5300 1.9550 ;
      RECT 0.0800 0.6700 1.5650 0.7600 ;
      RECT 1.4600 0.7600 1.5650 0.7800 ;
      RECT 1.4750 0.4100 1.5650 0.6700 ;
      RECT 1.9200 1.7550 2.0100 1.9900 ;
      RECT 1.9200 1.6200 2.0100 1.6650 ;
      RECT 0.0800 1.6650 2.3450 1.7550 ;
      RECT 2.2550 1.1800 2.3450 1.6650 ;
  END
END AND3_X4M_A12TH

MACRO AND3_X6M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.4450 0.3200 ;
        RECT 0.7050 0.3200 0.8750 0.5200 ;
        RECT 2.0550 0.3200 2.2250 0.5200 ;
        RECT 3.6700 0.3200 3.7600 0.5600 ;
        RECT 4.1900 0.3200 4.2800 0.6450 ;
        RECT 4.7100 0.3200 4.8000 0.6450 ;
        RECT 5.2300 0.3200 5.3200 0.6450 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.4450 2.7200 ;
        RECT 1.5750 1.8250 1.6650 2.0800 ;
        RECT 2.0950 1.8250 2.1850 2.0800 ;
        RECT 2.6150 1.8250 2.7050 2.0800 ;
        RECT 3.1350 1.8250 3.2250 2.0800 ;
        RECT 3.6700 1.8250 3.7600 2.0800 ;
        RECT 4.1900 1.7700 4.2800 2.0800 ;
        RECT 4.7100 1.7700 4.8000 2.0800 ;
        RECT 5.2300 1.7700 5.3200 2.0800 ;
    END
  END VDD

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 0.9200 3.5900 1.2050 ;
        RECT 0.7900 0.8300 3.5900 0.9200 ;
        RECT 0.7900 0.9200 0.8800 1.0250 ;
        RECT 2.0400 0.9200 2.2400 1.0750 ;
        RECT 0.5750 1.0250 0.8800 1.1150 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3750 1.4650 3.3300 1.5550 ;
        RECT 0.3750 1.4500 1.0600 1.4650 ;
        RECT 1.6500 1.4500 2.6200 1.4650 ;
        RECT 3.2400 1.2350 3.3300 1.4650 ;
        RECT 0.3750 1.1750 0.4650 1.4500 ;
        RECT 0.9700 1.1150 1.0600 1.4500 ;
        RECT 1.6500 1.3450 1.8750 1.4500 ;
        RECT 2.5300 1.2550 2.6200 1.4500 ;
        RECT 0.9700 1.0250 1.2100 1.1150 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1700 1.2500 1.5400 1.3750 ;
        RECT 1.4500 1.1200 1.5400 1.2500 ;
        RECT 1.4500 1.0300 1.9500 1.1200 ;
        RECT 1.8600 1.1200 1.9500 1.1650 ;
        RECT 1.8600 1.1650 2.4200 1.2550 ;
        RECT 2.3300 1.0750 3.1000 1.1650 ;
    END
    ANTENNAGATEAREA 0.3288 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.9450 5.1500 1.4500 ;
        RECT 3.9250 1.4500 5.1500 1.5500 ;
        RECT 3.9250 0.8450 5.1500 0.9450 ;
        RECT 3.9250 1.5500 4.0250 1.8850 ;
        RECT 4.4450 1.5500 4.5450 1.8850 ;
        RECT 4.9650 1.5500 5.0650 1.8850 ;
        RECT 3.9250 0.5000 4.0250 0.8450 ;
        RECT 4.4450 0.5000 4.5450 0.8450 ;
        RECT 4.9650 0.5000 5.0650 0.8450 ;
    END
    ANTENNADIFFAREA 0.975 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 3.6800 1.0700 4.9350 1.1600 ;
      RECT 0.0800 0.7400 0.1700 1.6450 ;
      RECT 0.0800 0.4850 0.1700 0.6500 ;
      RECT 1.2750 1.7350 1.4450 1.9350 ;
      RECT 0.0800 0.6500 1.5450 0.7400 ;
      RECT 1.3750 0.4500 1.5450 0.6500 ;
      RECT 1.7950 1.7350 1.9650 1.9350 ;
      RECT 2.3150 1.7350 2.4850 1.9350 ;
      RECT 2.8350 1.7350 3.0050 1.9350 ;
      RECT 2.8350 0.4500 3.0050 0.6500 ;
      RECT 3.3550 1.7350 3.5250 1.9350 ;
      RECT 0.0800 1.6450 3.7700 1.7350 ;
      RECT 3.6800 1.1600 3.7700 1.6450 ;
      RECT 3.6800 0.7400 3.7700 1.0700 ;
      RECT 2.8350 0.6500 3.7700 0.7400 ;
  END
END AND3_X6M_A12TH

MACRO AND3_X8M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0800 0.3200 0.1700 0.6000 ;
        RECT 1.3750 0.3200 1.5450 0.5250 ;
        RECT 2.7350 0.3200 2.9050 0.5250 ;
        RECT 4.2650 0.3200 4.4350 0.5250 ;
        RECT 4.8700 0.3200 4.9600 0.6850 ;
        RECT 5.3900 0.3200 5.4800 0.6850 ;
        RECT 5.9100 0.3200 6.0000 0.6850 ;
        RECT 6.4300 0.3200 6.5200 0.6850 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 2.2550 1.8200 2.3450 2.0800 ;
        RECT 2.7750 1.8200 2.8650 2.0800 ;
        RECT 3.2950 1.8200 3.3850 2.0800 ;
        RECT 3.8150 1.8200 3.9050 2.0800 ;
        RECT 4.3500 1.8200 4.4400 2.0800 ;
        RECT 4.8700 1.7700 4.9600 2.0800 ;
        RECT 5.3900 1.7700 5.4800 2.0800 ;
        RECT 5.9100 1.7700 6.0000 2.0800 ;
        RECT 6.4300 1.7700 6.5200 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4100 1.2500 3.1900 1.3500 ;
        RECT 2.4100 1.2200 2.5300 1.2500 ;
        RECT 3.1000 1.2200 3.1900 1.2500 ;
        RECT 2.3500 1.0650 2.5300 1.2200 ;
        RECT 3.1000 1.0650 3.3100 1.2200 ;
        RECT 1.6350 0.9750 2.5300 1.0650 ;
        RECT 3.1000 0.9750 4.0600 1.0650 ;
        RECT 1.6350 1.0650 1.7250 1.3700 ;
        RECT 3.9700 1.0650 4.0600 1.2500 ;
        RECT 1.5150 1.3700 1.7250 1.4600 ;
    END
    ANTENNAGATEAREA 0.423 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.8850 2.7500 1.0700 ;
        RECT 1.4550 0.7950 2.7500 0.8850 ;
        RECT 2.6400 1.0700 3.0100 1.1600 ;
        RECT 1.4550 0.8850 1.5450 1.1100 ;
        RECT 2.9200 0.8850 3.0100 1.0700 ;
        RECT 0.1850 1.1100 1.5450 1.2000 ;
        RECT 2.9200 0.7950 4.2900 0.8850 ;
        RECT 0.1850 1.2000 0.2750 1.3200 ;
        RECT 4.2000 0.8850 4.2900 1.2500 ;
    END
    ANTENNAGATEAREA 0.423 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6100 1.4500 0.9800 1.5500 ;
        RECT 0.6100 1.5500 1.9050 1.6400 ;
        RECT 1.8150 1.2450 1.9050 1.5500 ;
        RECT 1.8150 1.1550 2.2600 1.2450 ;
        RECT 2.1700 1.2450 2.2600 1.4400 ;
        RECT 2.1700 1.4400 3.5000 1.5300 ;
        RECT 3.4100 1.2550 3.5000 1.4400 ;
        RECT 3.4100 1.1550 3.8100 1.2550 ;
    END
    ANTENNAGATEAREA 0.423 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0350 0.9650 6.1650 1.4350 ;
        RECT 4.5900 1.4350 6.1650 1.4400 ;
        RECT 4.5900 0.9500 6.1650 0.9650 ;
        RECT 4.5900 1.4400 6.2800 1.5650 ;
        RECT 4.5900 0.8350 6.2800 0.9500 ;
        RECT 4.5900 1.5650 4.7200 1.8450 ;
        RECT 5.1100 1.5650 5.2400 1.8450 ;
        RECT 5.6300 1.5650 5.7600 1.8450 ;
        RECT 6.1500 1.5650 6.2800 1.8450 ;
        RECT 4.5900 0.5550 4.7200 0.8350 ;
        RECT 5.1100 0.5550 5.2400 0.8350 ;
        RECT 5.6300 0.5550 5.7600 0.8350 ;
        RECT 6.1500 0.5550 6.2800 0.8350 ;
    END
    ANTENNADIFFAREA 1.3 ;
  END Y
  OBS
    LAYER M1 ;
      RECT 4.3800 1.0850 5.9450 1.1750 ;
      RECT 0.7550 0.7050 0.8450 0.8350 ;
      RECT 0.7550 0.4650 0.8450 0.6150 ;
      RECT 1.9950 1.7100 2.0850 1.9900 ;
      RECT 2.0350 0.4150 2.2050 0.6150 ;
      RECT 2.5150 1.7100 2.6050 1.9900 ;
      RECT 3.0350 1.7100 3.1250 1.9900 ;
      RECT 3.5550 1.7100 3.6450 1.9900 ;
      RECT 3.5150 0.4150 3.6850 0.6150 ;
      RECT 4.0750 1.7100 4.1650 1.9900 ;
      RECT 1.9950 1.6200 4.4700 1.7100 ;
      RECT 4.3800 1.1750 4.4700 1.6200 ;
      RECT 4.3800 0.7050 4.4700 1.0850 ;
      RECT 0.7550 0.6150 4.4700 0.7050 ;
  END
END AND3_X8M_A12TH

MACRO AND4_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 1.6450 0.3200 ;
        RECT 1.0050 0.3200 1.1750 0.6700 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4500 0.8850 1.5500 1.5700 ;
        RECT 1.4050 1.5700 1.5500 1.6700 ;
        RECT 1.4050 0.7850 1.5500 0.8850 ;
        RECT 1.4050 1.6700 1.5050 1.9800 ;
        RECT 1.4050 0.4750 1.5050 0.7850 ;
    END
    ANTENNADIFFAREA 0.142625 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7000 1.0500 1.1100 1.1550 ;
    END
    ANTENNAGATEAREA 0.0459 ;
  END D

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9700 0.1600 1.3550 ;
    END
    ANTENNAGATEAREA 0.0459 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4400 1.0100 0.5600 1.3600 ;
    END
    ANTENNAGATEAREA 0.0459 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4950 1.4500 0.9150 1.5500 ;
    END
    ANTENNAGATEAREA 0.0459 ;
  END C

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 1.6450 2.7200 ;
        RECT 0.6100 1.8650 0.7100 2.0800 ;
        RECT 1.1450 1.8650 1.2450 2.0800 ;
        RECT 0.0900 1.8150 0.1900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.3550 1.6800 1.3000 1.7700 ;
      RECT 1.2100 1.2800 1.3000 1.6800 ;
      RECT 1.2100 1.1100 1.3450 1.2800 ;
      RECT 1.2100 0.8800 1.3000 1.1100 ;
      RECT 0.1300 0.7900 1.3000 0.8800 ;
      RECT 0.3550 1.7700 0.4450 1.9900 ;
      RECT 0.1300 0.4450 0.2200 0.7900 ;
      RECT 0.8750 1.7700 0.9650 1.9900 ;
  END
END AND4_X0P5M_A12TH

MACRO A2DFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.0000 3.5000 1.2000 ;
        RECT 3.4000 1.2000 3.5000 1.7100 ;
        RECT 3.4000 0.7100 3.5000 1.0000 ;
    END
    ANTENNADIFFAREA 0.1296 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0300 1.1450 4.1550 1.5000 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9700 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 0.3000 1.7300 0.4700 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9200 0.1750 1.3900 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7150 ;
        RECT 3.9150 0.3200 4.0850 0.8000 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5150 0.6950 1.6050 ;
      RECT 0.6050 1.6050 0.6950 1.7450 ;
      RECT 0.2650 0.7700 0.6450 0.8600 ;
      RECT 0.5550 0.6700 0.6450 0.7700 ;
      RECT 0.2650 0.8600 0.3550 1.5150 ;
      RECT 0.0800 1.6050 0.1700 1.7500 ;
      RECT 0.8000 1.6000 1.0300 1.6900 ;
      RECT 0.9300 1.0500 1.0300 1.6000 ;
      RECT 0.9300 0.9600 1.6400 1.0500 ;
      RECT 1.5500 1.0500 1.6400 1.2400 ;
      RECT 0.9300 0.6900 1.0200 0.9600 ;
      RECT 1.2300 1.6100 1.8400 1.7000 ;
      RECT 1.2300 1.1600 1.3200 1.6100 ;
      RECT 1.7500 0.6800 1.8400 1.6100 ;
      RECT 2.4400 1.3200 2.9500 1.4100 ;
      RECT 2.4400 0.9700 2.5400 1.3200 ;
      RECT 2.8600 0.9400 2.9500 1.3200 ;
      RECT 2.7800 0.8500 2.9500 0.9400 ;
      RECT 2.0100 0.7600 2.1000 1.7250 ;
      RECT 2.0100 0.6700 3.1500 0.7600 ;
      RECT 3.0600 0.7600 3.1500 1.2600 ;
      RECT 3.6100 1.6400 3.8100 1.7300 ;
      RECT 3.6100 0.8200 3.7000 1.6400 ;
      RECT 3.6100 0.7200 3.8050 0.8200 ;
      RECT 3.6100 0.5700 3.7050 0.7200 ;
      RECT 0.7400 0.4800 3.7050 0.5700 ;
      RECT 0.7400 0.5700 0.8300 1.4300 ;
      RECT 1.8800 0.4150 2.0850 0.4800 ;
      RECT 0.9300 1.8300 4.2150 1.9200 ;
      RECT 4.1250 1.7700 4.2150 1.8300 ;
      RECT 4.1250 1.6000 4.3350 1.7700 ;
      RECT 4.2450 1.0250 4.3350 1.6000 ;
      RECT 3.8250 0.9350 4.3350 1.0250 ;
      RECT 4.2300 0.6650 4.3350 0.9350 ;
      RECT 2.2150 0.9400 2.3050 1.8300 ;
  END
END A2DFFQN_X0P5M_A12TH

MACRO A2DFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6650 ;
        RECT 3.0550 0.3200 3.2250 0.3600 ;
        RECT 3.8950 0.3200 4.0650 0.7900 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2500 1.0100 3.4750 1.1900 ;
        RECT 3.3850 1.1900 3.4750 1.7100 ;
        RECT 3.3850 0.7300 3.4750 1.0100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8100 1.2500 4.1300 1.3500 ;
        RECT 4.0250 1.1350 4.1300 1.2500 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9600 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 1.4200 1.9500 1.5300 2.0800 ;
        RECT 2.6150 1.8950 2.7350 2.0800 ;
        RECT 0.3000 1.7100 0.4700 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9200 0.1750 1.3900 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5150 0.6950 1.6050 ;
      RECT 0.6050 1.6050 0.6950 1.7250 ;
      RECT 0.2650 0.7200 0.6450 0.8100 ;
      RECT 0.5550 0.5850 0.6450 0.7200 ;
      RECT 0.2650 0.8100 0.3550 1.5150 ;
      RECT 0.0800 1.6050 0.1700 1.7450 ;
      RECT 0.8000 1.5400 1.0300 1.6300 ;
      RECT 0.9300 1.0400 1.0300 1.5400 ;
      RECT 0.9300 0.9500 1.6400 1.0400 ;
      RECT 1.5500 1.0400 1.6400 1.2350 ;
      RECT 0.9300 0.6800 1.0200 0.9500 ;
      RECT 1.2350 1.5100 1.8450 1.6000 ;
      RECT 1.2350 1.1600 1.3250 1.5100 ;
      RECT 1.7550 0.6600 1.8450 1.5100 ;
      RECT 2.4650 1.3200 2.9700 1.4100 ;
      RECT 2.4650 0.9700 2.5550 1.3200 ;
      RECT 2.8800 0.9400 2.9700 1.3200 ;
      RECT 2.8000 0.8500 2.9700 0.9400 ;
      RECT 1.9350 1.5100 2.1100 1.6000 ;
      RECT 2.0200 0.7600 2.1100 1.5100 ;
      RECT 2.0200 0.6700 3.1600 0.7600 ;
      RECT 3.0700 0.7600 3.1600 1.2100 ;
      RECT 3.5950 1.5150 3.7900 1.6050 ;
      RECT 3.5950 0.8000 3.6850 1.5150 ;
      RECT 3.5950 0.7000 3.7850 0.8000 ;
      RECT 3.5950 0.5700 3.6850 0.7000 ;
      RECT 0.7400 0.4800 3.6850 0.5700 ;
      RECT 0.7400 0.5700 0.8300 1.4300 ;
      RECT 1.9000 0.4100 2.0850 0.4800 ;
      RECT 3.0300 1.8150 4.1950 1.9150 ;
      RECT 4.1050 1.6450 4.1950 1.8150 ;
      RECT 4.1050 1.4750 4.3100 1.6450 ;
      RECT 4.2200 1.0250 4.3100 1.4750 ;
      RECT 3.8050 0.9350 4.3100 1.0250 ;
      RECT 4.2100 0.6250 4.3100 0.9350 ;
      RECT 1.2100 1.7150 3.1200 1.8000 ;
      RECT 1.8500 1.8000 3.1200 1.8050 ;
      RECT 3.0300 1.8050 3.1200 1.8150 ;
      RECT 0.9100 1.8800 1.3000 1.9700 ;
      RECT 1.2100 1.8000 1.3000 1.8800 ;
      RECT 1.2100 1.7100 2.3100 1.7150 ;
      RECT 1.8500 1.8050 2.0200 1.9200 ;
      RECT 2.2200 0.8700 2.3100 1.7100 ;
  END
END A2DFFQN_X1M_A12TH

MACRO A2DFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.6450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6400 ;
        RECT 3.0550 0.3200 3.2250 0.3600 ;
        RECT 3.6100 0.3200 4.0000 0.3600 ;
        RECT 4.1150 0.3200 4.2850 0.7250 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3900 1.2500 3.7000 1.3500 ;
        RECT 3.3900 1.3500 3.4800 1.7100 ;
        RECT 3.6000 0.9500 3.7000 1.2500 ;
        RECT 3.3800 0.8500 3.7000 0.9500 ;
        RECT 3.3800 0.7050 3.4800 0.8500 ;
    END
    ANTENNADIFFAREA 0.328575 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0050 1.2500 4.3500 1.3500 ;
        RECT 4.2450 1.1350 4.3500 1.2500 ;
    END
    ANTENNAGATEAREA 0.0354 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 0.9600 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.6450 2.7200 ;
        RECT 1.4200 1.9500 1.5300 2.0800 ;
        RECT 2.6150 1.8650 2.7350 2.0800 ;
        RECT 0.3350 1.7550 0.4350 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9200 0.1750 1.3900 ;
    END
    ANTENNAGATEAREA 0.0672 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5150 0.6950 1.6050 ;
      RECT 0.6050 1.6050 0.6950 1.7900 ;
      RECT 0.2650 0.6100 0.6450 0.7000 ;
      RECT 0.5550 0.4750 0.6450 0.6100 ;
      RECT 0.2650 0.7000 0.3550 1.5150 ;
      RECT 0.0800 1.6050 0.1700 1.9250 ;
      RECT 0.8000 1.5400 1.0400 1.6300 ;
      RECT 0.9400 1.0400 1.0400 1.5400 ;
      RECT 0.9400 0.9500 1.6250 1.0400 ;
      RECT 1.5350 1.0400 1.6250 1.2350 ;
      RECT 0.9400 0.6800 1.0300 0.9500 ;
      RECT 1.2450 1.5000 1.8450 1.5900 ;
      RECT 1.2450 1.1600 1.3350 1.5000 ;
      RECT 1.7550 0.7300 1.8450 1.5000 ;
      RECT 2.4650 1.3200 2.8850 1.4100 ;
      RECT 2.4650 0.9700 2.5550 1.3200 ;
      RECT 2.7950 0.9450 2.8850 1.3200 ;
      RECT 2.7950 0.8500 2.9700 0.9450 ;
      RECT 3.0850 1.0600 3.4900 1.1500 ;
      RECT 1.9350 1.4550 2.1100 1.5450 ;
      RECT 2.0200 0.7600 2.1100 1.4550 ;
      RECT 2.0200 0.6700 3.1750 0.7600 ;
      RECT 3.0850 0.7600 3.1750 1.0600 ;
      RECT 3.8100 1.5150 4.0100 1.6050 ;
      RECT 3.8100 0.6750 4.0050 0.7750 ;
      RECT 3.8100 0.7750 3.9000 1.5150 ;
      RECT 3.8100 0.5700 3.9050 0.6750 ;
      RECT 0.7400 0.4800 3.9050 0.5700 ;
      RECT 0.7400 0.5700 0.8300 1.4300 ;
      RECT 1.9000 0.4150 2.0900 0.4800 ;
      RECT 3.0300 1.8150 4.4150 1.9150 ;
      RECT 4.3250 1.6450 4.4150 1.8150 ;
      RECT 4.3250 1.4750 4.5300 1.6450 ;
      RECT 4.4400 1.0250 4.5300 1.4750 ;
      RECT 4.0250 0.9350 4.5300 1.0250 ;
      RECT 4.4300 0.6250 4.5300 0.9350 ;
      RECT 1.2100 1.6850 3.1200 1.7700 ;
      RECT 1.8500 1.7700 3.1200 1.7750 ;
      RECT 3.0300 1.7750 3.1200 1.8150 ;
      RECT 0.9550 1.8800 1.3000 1.9700 ;
      RECT 1.2100 1.7700 1.3000 1.8800 ;
      RECT 1.2100 1.6800 2.3100 1.6850 ;
      RECT 1.8500 1.7750 2.0200 1.9900 ;
      RECT 2.2200 0.8700 2.3100 1.6800 ;
  END
END A2DFFQN_X2M_A12TH

MACRO A2DFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.0950 0.3200 0.1950 0.6450 ;
        RECT 2.6050 0.3200 2.8150 0.3800 ;
        RECT 3.1100 0.3200 3.2800 0.3600 ;
        RECT 3.6600 0.3200 3.8300 0.3600 ;
        RECT 4.5150 0.3200 4.6350 0.6950 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3800 1.4500 4.0600 1.5500 ;
        RECT 3.9700 0.8200 4.0600 1.4500 ;
        RECT 3.3800 0.7300 4.0600 0.8200 ;
    END
    ANTENNADIFFAREA 0.593125 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6500 1.0100 4.7500 1.4300 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6100 1.2900 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 4.5200 1.8950 4.6300 2.0800 ;
        RECT 2.5500 1.8650 2.6700 2.0800 ;
        RECT 0.3550 1.7000 0.4550 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 1.0450 0.1750 1.3900 ;
    END
    ANTENNAGATEAREA 0.0798 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.1000 1.5100 0.7100 1.6000 ;
      RECT 0.6200 1.6000 0.7100 1.9200 ;
      RECT 0.2650 0.7750 0.6650 0.8650 ;
      RECT 0.5750 0.4350 0.6650 0.7750 ;
      RECT 0.2650 0.8650 0.3550 1.5100 ;
      RECT 0.1000 1.6000 0.1900 1.9200 ;
      RECT 0.8200 1.5300 1.0600 1.6200 ;
      RECT 0.9600 1.0400 1.0600 1.5300 ;
      RECT 0.9600 0.9500 1.6150 1.0400 ;
      RECT 1.5250 1.0400 1.6150 1.2350 ;
      RECT 0.9600 0.6800 1.0500 0.9500 ;
      RECT 1.2550 1.5000 1.8100 1.5900 ;
      RECT 1.2550 1.1600 1.3450 1.5000 ;
      RECT 1.7200 0.9050 1.8100 1.5000 ;
      RECT 1.7200 0.8150 1.9250 0.9050 ;
      RECT 2.4850 1.3800 2.9850 1.4700 ;
      RECT 2.4850 1.1500 2.5750 1.3800 ;
      RECT 2.8950 0.9450 2.9850 1.3800 ;
      RECT 2.8550 0.8500 3.0450 0.9450 ;
      RECT 3.1600 1.0850 3.5750 1.1750 ;
      RECT 1.9200 1.4800 2.1250 1.5700 ;
      RECT 2.0350 0.7600 2.1250 1.4800 ;
      RECT 2.0350 0.6700 3.2500 0.7600 ;
      RECT 3.1600 0.7600 3.2500 1.0850 ;
      RECT 4.2050 1.4200 4.3750 1.5300 ;
      RECT 4.2050 0.6050 4.2950 1.4200 ;
      RECT 4.2050 0.5700 4.3750 0.6050 ;
      RECT 0.7600 0.4800 4.3750 0.5700 ;
      RECT 0.7600 0.5700 0.8500 1.4300 ;
      RECT 2.2350 0.4100 2.4100 0.4800 ;
      RECT 0.9500 1.8600 1.2250 1.9500 ;
      RECT 1.1350 1.7700 1.2250 1.8600 ;
      RECT 1.1350 1.6850 4.5900 1.7700 ;
      RECT 1.1350 1.6800 2.3250 1.6850 ;
      RECT 2.1250 1.7700 4.5900 1.7750 ;
      RECT 2.2350 1.0000 2.3250 1.6800 ;
      RECT 4.3900 0.8300 4.9500 0.9200 ;
      RECT 4.5000 1.5400 4.9500 1.6300 ;
      RECT 4.5000 1.6300 4.5900 1.6850 ;
      RECT 4.7550 0.6000 4.9500 0.6900 ;
      RECT 4.8600 0.6900 4.9500 0.8300 ;
      RECT 4.8600 0.9200 4.9500 1.5400 ;
      RECT 2.1250 1.6850 2.3500 1.9600 ;
      RECT 2.1250 1.6800 2.3250 1.6850 ;
  END
END A2DFFQN_X3M_A12TH

MACRO A2DFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.7000 ;
        RECT 1.4850 0.3200 1.5850 0.8450 ;
        RECT 2.6050 0.3200 2.7050 0.8450 ;
        RECT 3.1150 0.3200 3.2150 0.9900 ;
        RECT 3.9000 0.3200 4.0000 0.8900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5250 1.8500 0.8150 1.9500 ;
        RECT 0.5250 1.6500 0.6250 1.8500 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.0550 3.5500 1.6500 ;
        RECT 3.3050 1.6500 3.5500 1.7400 ;
        RECT 3.3750 0.9550 3.5500 1.0550 ;
        RECT 3.3750 0.7550 3.4750 0.9550 ;
    END
    ANTENNADIFFAREA 0.14175 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0100 0.9900 4.1500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0207 ;
  END CK

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 0.8500 0.3900 1.0050 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 2.4850 1.8700 2.5850 2.0800 ;
        RECT 4.0200 1.8400 4.1900 2.0800 ;
        RECT 0.3350 1.3400 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5450 1.3750 0.7300 1.4650 ;
      RECT 0.5450 1.2500 0.6350 1.3750 ;
      RECT 0.0800 1.1600 0.6350 1.2500 ;
      RECT 0.5450 0.8150 0.6350 1.1600 ;
      RECT 0.5450 0.7250 0.6900 0.8150 ;
      RECT 0.6000 0.6050 0.6900 0.7250 ;
      RECT 0.0800 1.2500 0.1700 1.5400 ;
      RECT 0.7250 1.0600 0.8700 1.2500 ;
      RECT 0.7800 0.5450 0.8700 1.0600 ;
      RECT 0.7800 0.4550 1.2000 0.5450 ;
      RECT 0.8200 1.3950 1.6550 1.4850 ;
      RECT 1.5650 1.2750 1.6550 1.3950 ;
      RECT 0.8200 1.3900 1.1300 1.3950 ;
      RECT 1.0400 0.6350 1.1300 1.3900 ;
      RECT 1.6450 1.6250 1.8400 1.7150 ;
      RECT 1.7500 1.0950 1.8400 1.6250 ;
      RECT 1.3250 1.0050 1.8400 1.0950 ;
      RECT 1.7500 0.6350 1.8400 1.0050 ;
      RECT 2.7050 1.0550 2.7950 1.2700 ;
      RECT 2.4250 0.9650 2.7950 1.0550 ;
      RECT 2.4250 0.7850 2.5150 0.9650 ;
      RECT 1.9700 0.6950 2.5150 0.7850 ;
      RECT 1.9700 0.7850 2.0600 1.7400 ;
      RECT 2.8750 1.5350 3.3050 1.5600 ;
      RECT 2.4100 1.4450 3.3050 1.5350 ;
      RECT 3.2150 1.1500 3.3050 1.4450 ;
      RECT 2.4100 1.1650 2.5000 1.4450 ;
      RECT 2.8750 1.5600 2.9650 1.7400 ;
      RECT 2.9350 0.7850 3.0250 1.4450 ;
      RECT 2.8150 0.6950 3.0250 0.7850 ;
      RECT 3.6400 0.5050 3.7300 1.5250 ;
      RECT 3.4500 0.4150 3.7300 0.5050 ;
      RECT 3.8250 1.5100 4.3500 1.6000 ;
      RECT 4.2250 1.3600 4.3500 1.5100 ;
      RECT 4.2600 0.8850 4.3500 1.3600 ;
      RECT 4.1900 0.6800 4.3500 0.8850 ;
      RECT 2.6750 1.8300 3.9150 1.9200 ;
      RECT 3.8250 1.6000 3.9150 1.8300 ;
      RECT 3.8250 1.0100 3.9150 1.5100 ;
      RECT 1.8200 1.9200 1.9900 1.9650 ;
      RECT 0.9900 1.8300 2.2650 1.9200 ;
      RECT 2.1750 1.7350 2.2650 1.8300 ;
      RECT 2.1750 0.9050 2.2650 1.6450 ;
      RECT 2.1750 1.6450 2.7650 1.7350 ;
      RECT 2.6750 1.7350 2.7650 1.8300 ;
  END
END A2DFFQ_X0P5M_A12TH

MACRO A2DFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.4450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.6200 ;
        RECT 1.4850 0.3200 1.5850 0.8450 ;
        RECT 2.6050 0.3200 2.7050 0.8450 ;
        RECT 3.9000 0.3200 4.0000 0.8900 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5250 1.8500 0.8150 1.9500 ;
        RECT 0.5250 1.6500 0.6250 1.8500 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END A

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4500 1.0550 3.5500 1.6500 ;
        RECT 3.3050 1.6500 3.5500 1.7400 ;
        RECT 3.3750 0.9550 3.5500 1.0550 ;
        RECT 3.3750 0.7150 3.4750 0.9550 ;
    END
    ANTENNADIFFAREA 0.266075 ;
  END Q

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0100 0.9900 4.1500 1.3000 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END CK

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1000 0.8500 0.3900 1.0050 ;
    END
    ANTENNAGATEAREA 0.0408 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.4450 2.7200 ;
        RECT 4.0200 1.8400 4.1900 2.0800 ;
        RECT 2.4850 1.8300 2.5850 2.0800 ;
        RECT 0.3350 1.4250 0.4350 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5450 1.3750 0.7300 1.4650 ;
      RECT 0.5450 1.2500 0.6350 1.3750 ;
      RECT 0.0800 1.1600 0.6350 1.2500 ;
      RECT 0.5450 0.8150 0.6350 1.1600 ;
      RECT 0.5450 0.7250 0.6900 0.8150 ;
      RECT 0.6000 0.6050 0.6900 0.7250 ;
      RECT 0.0800 1.2500 0.1700 1.5700 ;
      RECT 0.7250 1.0600 0.8700 1.2500 ;
      RECT 0.7800 0.5450 0.8700 1.0600 ;
      RECT 0.7800 0.4550 1.2000 0.5450 ;
      RECT 0.8200 1.3950 1.6550 1.4850 ;
      RECT 1.5650 1.2750 1.6550 1.3950 ;
      RECT 0.8200 1.3900 1.1150 1.3950 ;
      RECT 1.0250 0.6350 1.1150 1.3900 ;
      RECT 1.6100 1.6250 1.8400 1.7150 ;
      RECT 1.7500 1.0950 1.8400 1.6250 ;
      RECT 1.3250 1.0050 1.8400 1.0950 ;
      RECT 1.7500 0.6350 1.8400 1.0050 ;
      RECT 2.7050 1.0550 2.7950 1.2700 ;
      RECT 2.4250 0.9650 2.7950 1.0550 ;
      RECT 2.4250 0.7850 2.5150 0.9650 ;
      RECT 1.9650 0.6950 2.5150 0.7850 ;
      RECT 1.9650 0.7850 2.0550 1.7400 ;
      RECT 2.8750 1.5600 2.9650 1.7200 ;
      RECT 2.8750 1.5350 3.0250 1.5600 ;
      RECT 2.4100 1.4450 3.0250 1.5350 ;
      RECT 2.9350 1.1650 3.0250 1.4450 ;
      RECT 2.9350 1.0750 3.2650 1.1650 ;
      RECT 2.9350 0.7850 3.0250 1.0750 ;
      RECT 2.8150 0.6950 3.0250 0.7850 ;
      RECT 2.4100 1.1650 2.5000 1.4450 ;
      RECT 3.6400 0.5850 3.7300 1.5250 ;
      RECT 3.1300 0.5000 3.7300 0.5850 ;
      RECT 2.8950 0.4950 3.7300 0.5000 ;
      RECT 2.8950 0.4100 3.2200 0.4950 ;
      RECT 3.8250 1.5100 4.3500 1.6000 ;
      RECT 4.2250 1.3600 4.3500 1.5100 ;
      RECT 4.2600 0.8850 4.3500 1.3600 ;
      RECT 4.1900 0.6800 4.3500 0.8850 ;
      RECT 2.6950 1.8300 3.9150 1.9200 ;
      RECT 3.8250 1.6000 3.9150 1.8300 ;
      RECT 3.8250 1.0100 3.9150 1.5100 ;
      RECT 1.8150 1.9200 1.9850 1.9900 ;
      RECT 0.9900 1.8300 2.2650 1.9200 ;
      RECT 2.1750 1.7350 2.2650 1.8300 ;
      RECT 2.1750 0.9050 2.2650 1.6450 ;
      RECT 2.1750 1.6450 2.7850 1.7350 ;
      RECT 2.6950 1.7350 2.7850 1.8300 ;
  END
END A2DFFQ_X1M_A12TH

MACRO A2DFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.8450 0.3200 ;
        RECT 0.0750 0.3200 0.1750 0.8800 ;
        RECT 1.4400 0.3200 1.5400 0.7600 ;
        RECT 3.2500 0.3200 3.3500 0.4600 ;
        RECT 3.7750 0.3200 3.8750 0.4600 ;
        RECT 4.3250 0.3200 4.4250 0.8900 ;
    END
  END VSS

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0450 1.0250 0.1600 1.4100 ;
    END
    ANTENNAGATEAREA 0.0528 ;
  END B

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8500 0.9000 3.9500 1.3600 ;
        RECT 3.4600 1.3600 3.9500 1.4600 ;
        RECT 3.4600 0.8000 3.9500 0.9000 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.8450 2.7200 ;
        RECT 1.3550 1.9150 1.5350 2.0800 ;
        RECT 2.6950 1.8200 2.7950 2.0800 ;
        RECT 3.2450 1.8000 3.3450 2.0800 ;
        RECT 3.7750 1.8000 3.8750 2.0800 ;
        RECT 4.3300 1.8000 4.4200 2.0800 ;
        RECT 0.3350 1.7050 0.4350 2.0800 ;
    END
  END VDD

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4150 1.0100 4.5550 1.3450 ;
    END
    ANTENNAGATEAREA 0.0291 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.9800 0.5500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0528 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0800 1.5000 0.6900 1.5900 ;
      RECT 0.6000 1.5900 0.6900 1.8900 ;
      RECT 0.2650 0.7800 0.6300 0.8700 ;
      RECT 0.5400 0.4600 0.6300 0.7800 ;
      RECT 0.2650 0.8700 0.3550 1.5000 ;
      RECT 0.0800 1.5900 0.1700 1.8900 ;
      RECT 0.6600 1.2950 0.8500 1.3850 ;
      RECT 0.7600 0.5450 0.8500 1.2950 ;
      RECT 0.7600 0.4550 1.1800 0.5450 ;
      RECT 0.9400 1.0500 1.6500 1.1400 ;
      RECT 1.5600 1.1400 1.6500 1.2600 ;
      RECT 0.8000 1.5300 1.0400 1.6200 ;
      RECT 0.9400 1.1400 1.0400 1.5300 ;
      RECT 0.9400 0.6550 1.0300 1.0500 ;
      RECT 1.2450 1.4650 1.8400 1.5550 ;
      RECT 1.2450 1.2350 1.3350 1.4650 ;
      RECT 1.7500 1.1850 1.8400 1.4650 ;
      RECT 1.7500 1.0950 1.8900 1.1850 ;
      RECT 1.8000 0.8150 1.8900 1.0950 ;
      RECT 1.9300 1.4050 2.0950 1.5900 ;
      RECT 2.0050 0.7500 2.0950 1.4050 ;
      RECT 2.0050 0.6600 2.8100 0.7500 ;
      RECT 2.7200 0.7500 2.8100 1.0100 ;
      RECT 2.7200 1.0100 2.9000 1.1000 ;
      RECT 2.8100 1.1000 2.9000 1.2200 ;
      RECT 3.0250 1.0850 3.7550 1.1750 ;
      RECT 2.4750 1.4200 3.1150 1.5100 ;
      RECT 3.0250 1.1750 3.1150 1.4200 ;
      RECT 2.4750 1.0650 2.5650 1.4200 ;
      RECT 3.0250 0.8900 3.1150 1.0850 ;
      RECT 2.9050 0.8000 3.1150 0.8900 ;
      RECT 4.0450 0.6900 4.1350 1.4700 ;
      RECT 2.9650 0.6000 4.1350 0.6900 ;
      RECT 2.9650 0.5700 3.0550 0.6000 ;
      RECT 1.9150 0.4800 3.0550 0.5700 ;
      RECT 1.9150 0.4200 2.0850 0.4800 ;
      RECT 1.1150 1.6850 4.7450 1.7100 ;
      RECT 2.2350 1.6200 4.7450 1.6850 ;
      RECT 4.6100 1.4500 4.7450 1.6200 ;
      RECT 4.6550 0.8250 4.7450 1.4500 ;
      RECT 4.5550 0.7350 4.7450 0.8250 ;
      RECT 0.9400 1.8800 1.2050 1.9700 ;
      RECT 1.1150 1.7750 1.2050 1.8800 ;
      RECT 1.1150 1.7100 2.3250 1.7750 ;
      RECT 1.8300 1.7750 2.0000 1.9500 ;
      RECT 2.2350 0.8400 2.3250 1.6200 ;
      RECT 4.0950 1.7100 4.1900 1.8250 ;
      RECT 4.1000 1.8250 4.1900 1.9200 ;
  END
END A2DFFQ_X2M_A12TH

MACRO A2DFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.0450 0.3200 ;
        RECT 0.5300 0.3200 0.7000 0.3950 ;
        RECT 2.0500 0.3200 2.1500 0.8850 ;
        RECT 3.2500 0.3200 3.3500 0.7550 ;
        RECT 3.9750 0.3200 4.0750 0.4300 ;
        RECT 4.5650 0.3200 4.6650 0.6000 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.2200 4.1500 1.4100 ;
        RECT 3.9750 1.0500 4.1500 1.2200 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CK

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5300 1.0100 0.7550 1.1200 ;
        RECT 0.6450 1.1200 0.7550 1.3500 ;
        RECT 0.5300 0.9200 0.6400 1.0100 ;
    END
    ANTENNAGATEAREA 0.0624 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0500 0.9200 0.1600 1.4000 ;
    END
    ANTENNAGATEAREA 0.0624 ;
  END A

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3050 1.2500 4.9500 1.3500 ;
        RECT 4.3050 1.3500 4.4050 1.7200 ;
        RECT 4.8300 1.3500 4.9500 1.7350 ;
        RECT 4.8500 0.9500 4.9500 1.2500 ;
        RECT 4.4250 0.8500 4.9500 0.9500 ;
        RECT 4.4250 0.7800 4.5250 0.8500 ;
        RECT 4.8300 0.5200 4.9500 0.8500 ;
        RECT 4.3050 0.6900 4.5250 0.7800 ;
        RECT 4.3050 0.4100 4.4050 0.6900 ;
    END
    ANTENNADIFFAREA 0.585 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.0450 2.7200 ;
        RECT 0.6350 1.8200 0.7350 2.0800 ;
        RECT 4.0450 2.0500 4.6650 2.0800 ;
        RECT 0.0750 1.5600 0.1750 2.0800 ;
        RECT 4.0450 1.7900 4.1450 2.0500 ;
        RECT 4.5650 1.7700 4.6650 2.0500 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 1.1650 1.7300 1.2550 1.9300 ;
      RECT 0.3350 1.6400 1.2550 1.7300 ;
      RECT 1.1650 1.5400 1.2550 1.6400 ;
      RECT 0.4700 0.4950 1.2700 0.5850 ;
      RECT 1.1800 0.5850 1.2700 0.9150 ;
      RECT 0.3350 0.7800 0.4400 1.6400 ;
      RECT 0.0800 0.4100 0.1700 0.6900 ;
      RECT 0.0800 0.6900 0.5600 0.7800 ;
      RECT 0.4700 0.5850 0.5600 0.6900 ;
      RECT 0.9300 1.2450 1.0200 1.5350 ;
      RECT 0.9300 1.1550 1.5000 1.2450 ;
      RECT 0.9300 0.6750 1.0200 1.1550 ;
      RECT 1.6500 1.0200 2.2200 1.1100 ;
      RECT 1.4200 1.5650 1.7400 1.6550 ;
      RECT 1.6500 1.1100 1.7400 1.5650 ;
      RECT 1.6500 0.8550 1.7400 1.0200 ;
      RECT 1.4350 0.7650 1.7400 0.8550 ;
      RECT 1.8750 1.2350 2.4050 1.3250 ;
      RECT 2.3150 1.3250 2.4050 1.7200 ;
      RECT 2.3150 0.4700 2.4050 1.2350 ;
      RECT 1.8750 1.3250 1.9650 1.4350 ;
      RECT 2.9400 0.8900 3.4300 0.9800 ;
      RECT 2.7200 1.4400 2.8100 1.5500 ;
      RECT 2.7200 1.3500 3.0300 1.4400 ;
      RECT 2.9400 0.9800 3.0300 1.3500 ;
      RECT 2.9400 0.5700 3.0300 0.8900 ;
      RECT 2.6000 0.4800 3.0300 0.5700 ;
      RECT 1.6050 1.8200 3.8650 1.9100 ;
      RECT 3.7750 0.7900 3.8650 1.8200 ;
      RECT 2.5150 1.2600 2.6050 1.8200 ;
      RECT 2.5150 1.1700 2.8450 1.2600 ;
      RECT 2.7550 0.6900 2.8450 1.1700 ;
      RECT 4.2450 1.0600 4.6550 1.1500 ;
      RECT 3.5100 1.2600 3.6200 1.6700 ;
      RECT 3.1400 1.0900 3.6200 1.2600 ;
      RECT 3.5200 0.7000 3.6200 1.0900 ;
      RECT 3.5200 0.4100 3.6200 0.6100 ;
      RECT 3.5200 0.6100 4.0650 0.7000 ;
      RECT 3.9750 0.7000 4.0650 0.8700 ;
      RECT 3.9750 0.8700 4.3350 0.9600 ;
      RECT 4.2450 0.9600 4.3350 1.0600 ;
  END
END A2DFFQ_X3M_A12TH

MACRO A2DFFQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.5050 0.3200 0.6050 0.4300 ;
        RECT 1.0250 0.3200 1.1250 0.4300 ;
        RECT 1.5450 0.3200 1.6450 0.4200 ;
        RECT 2.9350 0.3200 3.0350 0.5000 ;
        RECT 4.2650 0.3200 4.3650 0.4400 ;
        RECT 5.0450 0.3200 5.1450 0.6500 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8550 1.4500 1.5500 1.5500 ;
        RECT 0.8550 1.5500 0.9550 1.8800 ;
        RECT 1.3750 1.5500 1.4750 1.8800 ;
        RECT 1.4500 0.8850 1.5500 1.4500 ;
        RECT 0.7100 0.7850 1.5500 0.8850 ;
    END
    ANTENNADIFFAREA 0.65 ;
  END Q

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3000 1.0500 4.7300 1.1500 ;
        RECT 4.6300 0.9550 4.7300 1.0500 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.7300 4.9600 1.1850 ;
    END
    ANTENNAGATEAREA 0.069 ;
  END B

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2100 1.0000 5.3500 1.3800 ;
    END
    ANTENNAGATEAREA 0.0381 ;
  END CK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.5950 1.7700 0.6950 2.0800 ;
        RECT 1.1150 2.0500 1.7350 2.0800 ;
        RECT 0.0750 1.7500 0.1750 2.0800 ;
        RECT 5.1350 1.7100 5.2350 2.0800 ;
        RECT 1.1150 1.7700 1.2150 2.0500 ;
        RECT 1.6350 1.7700 1.7350 2.0500 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.2250 1.0850 1.2800 1.1750 ;
      RECT 0.3400 1.6350 0.4300 1.9650 ;
      RECT 0.2250 0.7400 0.3150 1.0850 ;
      RECT 0.3400 1.5350 0.7550 1.6350 ;
      RECT 0.6650 1.1750 0.7550 1.5350 ;
      RECT 2.2100 1.5300 2.3000 1.8300 ;
      RECT 1.6600 1.4400 2.3000 1.5300 ;
      RECT 1.6600 0.6100 1.7500 1.4400 ;
      RECT 0.0450 0.5200 1.9100 0.6100 ;
      RECT 1.8100 0.4300 2.2250 0.5200 ;
      RECT 0.0450 0.6100 0.1350 1.3350 ;
      RECT 0.0450 1.3350 0.5750 1.4250 ;
      RECT 2.5700 1.5400 2.6600 1.6400 ;
      RECT 2.5700 1.4450 2.7750 1.5400 ;
      RECT 2.6850 0.9200 2.7750 1.4450 ;
      RECT 2.5050 0.8300 3.2450 0.9200 ;
      RECT 2.5050 0.6800 2.6050 0.8300 ;
      RECT 3.4750 1.2000 3.5650 1.6400 ;
      RECT 2.8650 1.1100 3.5650 1.2000 ;
      RECT 2.8650 1.0300 2.9550 1.1100 ;
      RECT 3.4700 0.7750 3.5650 1.1100 ;
      RECT 3.4700 0.6800 3.6550 0.7750 ;
      RECT 3.7450 1.6500 4.1550 1.7400 ;
      RECT 3.7450 0.5700 3.8350 1.6500 ;
      RECT 3.2600 0.4800 4.1400 0.5700 ;
      RECT 3.2600 0.5700 3.3500 0.6200 ;
      RECT 3.9700 0.4100 4.1400 0.4800 ;
      RECT 2.7500 0.6200 3.3500 0.7100 ;
      RECT 2.7500 0.5700 2.8400 0.6200 ;
      RECT 2.3150 0.4800 2.8400 0.5700 ;
      RECT 2.3150 0.5700 2.4050 0.9300 ;
      RECT 2.0350 0.9300 2.4050 1.0200 ;
      RECT 2.0450 1.0200 2.1350 1.1500 ;
      RECT 4.7400 1.5100 4.8300 1.6900 ;
      RECT 4.5100 1.4200 4.8300 1.5100 ;
      RECT 4.5100 1.3500 4.6000 1.4200 ;
      RECT 3.9300 1.2600 4.6000 1.3500 ;
      RECT 3.9300 0.6800 4.6100 0.7800 ;
      RECT 4.5200 0.4100 4.6100 0.6800 ;
      RECT 3.9300 1.3500 4.0250 1.5050 ;
      RECT 3.9300 0.7800 4.0250 1.2600 ;
      RECT 4.9200 1.5200 5.5450 1.6100 ;
      RECT 5.4100 1.6100 5.5450 1.9100 ;
      RECT 5.4450 0.7950 5.5450 1.5200 ;
      RECT 5.3600 0.6800 5.5450 0.7950 ;
      RECT 3.2700 1.8550 5.0100 1.9200 ;
      RECT 2.3900 1.8300 5.0100 1.8550 ;
      RECT 4.9200 1.6100 5.0100 1.8300 ;
      RECT 2.3900 1.7500 3.4450 1.8300 ;
      RECT 2.3900 1.3300 2.4800 1.7500 ;
      RECT 1.8450 1.2400 2.5950 1.3300 ;
      RECT 2.5050 1.0300 2.5950 1.2400 ;
      RECT 1.8450 0.8100 1.9350 1.2400 ;
      RECT 1.8450 0.7200 2.1000 0.8100 ;
      RECT 4.3050 1.5600 4.3950 1.8300 ;
      RECT 4.2050 1.4700 4.3950 1.5600 ;
  END
END A2DFFQ_X4M_A12TH

MACRO A2SDFFQN_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7400 ;
        RECT 0.9400 0.3200 1.1100 0.4350 ;
        RECT 2.6750 0.3200 2.8450 0.3900 ;
        RECT 3.8150 0.3200 3.9150 0.6750 ;
        RECT 5.1100 0.3200 5.2100 0.5750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.2100 5.0400 1.4800 ;
        RECT 4.9400 1.0750 5.0400 1.2100 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7800 4.5650 1.2900 ;
        RECT 4.3700 1.2900 4.5650 1.4700 ;
        RECT 4.3950 0.6800 4.5650 0.7800 ;
    END
    ANTENNADIFFAREA 0.153125 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.3100 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 1.0100 1.8300 1.1800 2.0800 ;
        RECT 0.3300 1.8050 0.4400 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.7900 1.8250 1.1600 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9000 1.5500 ;
        RECT 0.2500 1.5500 0.3600 1.6650 ;
        RECT 0.8000 1.0050 0.9000 1.4500 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.4400 1.5950 1.5500 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5700 1.2600 0.6600 ;
      RECT 1.1700 0.6600 1.2600 0.9000 ;
      RECT 0.0700 0.8300 0.7250 0.9200 ;
      RECT 0.6350 0.6600 0.7250 0.8300 ;
      RECT 0.0700 1.8050 0.2050 1.9750 ;
      RECT 0.0700 0.9200 0.1600 1.8050 ;
      RECT 0.0700 0.6850 0.1800 0.8300 ;
      RECT 1.2900 1.8300 2.0300 1.9200 ;
      RECT 0.8100 1.6500 1.9750 1.7400 ;
      RECT 1.8850 1.6100 1.9750 1.6500 ;
      RECT 1.8850 1.5200 2.0750 1.6100 ;
      RECT 1.3700 0.5200 1.9350 0.6100 ;
      RECT 1.8350 0.4200 1.9350 0.5200 ;
      RECT 0.9900 1.0100 1.4600 1.1000 ;
      RECT 1.3700 0.6100 1.4600 1.0100 ;
      RECT 0.9900 1.1000 1.0800 1.6500 ;
      RECT 0.9900 0.8500 1.0800 1.0100 ;
      RECT 0.8800 0.7500 1.0800 0.8500 ;
      RECT 0.8100 1.7400 0.9000 1.9900 ;
      RECT 2.2250 1.2400 2.3150 1.7400 ;
      RECT 2.2250 1.1400 2.9600 1.2400 ;
      RECT 2.8600 1.2400 2.9600 1.3500 ;
      RECT 2.2250 0.6800 2.3150 1.1400 ;
      RECT 3.0500 1.5950 3.2200 1.6950 ;
      RECT 3.0500 1.0500 3.1400 1.5950 ;
      RECT 2.5450 0.9600 3.1400 1.0500 ;
      RECT 3.0300 0.8150 3.1400 0.9600 ;
      RECT 3.0300 0.7150 3.2250 0.8150 ;
      RECT 3.3200 1.6050 4.0400 1.7050 ;
      RECT 3.9400 1.1850 4.0400 1.6050 ;
      RECT 3.3200 0.6800 3.4200 1.6050 ;
      RECT 3.6950 1.0750 3.7850 1.1800 ;
      RECT 3.6950 0.9850 4.2800 1.0750 ;
      RECT 4.1700 1.0750 4.2800 1.7350 ;
      RECT 4.1900 0.6800 4.2800 0.9850 ;
      RECT 2.4200 1.8300 5.3400 1.9200 ;
      RECT 5.2500 0.9750 5.3400 1.8300 ;
      RECT 4.7500 0.8850 5.3400 0.9750 ;
      RECT 4.7500 0.6800 4.8400 0.8850 ;
      RECT 2.4200 1.3500 2.5100 1.8300 ;
      RECT 4.9300 0.6850 5.5200 0.7750 ;
      RECT 5.4300 0.7750 5.5200 1.9650 ;
      RECT 1.9550 1.2900 2.1350 1.3800 ;
      RECT 2.0450 0.5700 2.1350 1.2900 ;
      RECT 2.0450 0.4800 3.6050 0.5700 ;
      RECT 3.5150 0.5700 3.6050 0.7850 ;
      RECT 3.5150 0.8750 3.6050 1.4900 ;
      RECT 4.0050 0.4800 5.0200 0.5700 ;
      RECT 4.9300 0.5700 5.0200 0.6850 ;
      RECT 3.5150 0.7850 4.0950 0.8750 ;
      RECT 4.0050 0.5700 4.0950 0.7850 ;
  END
END A2SDFFQN_X0P5M_A12TH

MACRO A2SDFFQN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7250 ;
        RECT 0.8850 0.3200 1.2550 0.3850 ;
        RECT 3.7900 0.3200 4.1600 0.3900 ;
        RECT 5.3400 0.3200 5.4500 0.6400 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 1.0100 5.6350 1.1900 ;
        RECT 5.5300 1.1900 5.6350 1.4150 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6200 0.6600 4.7500 1.7100 ;
    END
    ANTENNADIFFAREA 0.2448 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.2000 ;
        RECT 0.4500 1.2000 0.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 3.7900 2.0200 4.1600 2.0800 ;
        RECT 2.9150 1.9050 3.0850 2.0800 ;
        RECT 0.3350 1.6900 0.4450 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4850 1.0500 1.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.0666 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9000 1.5500 ;
        RECT 0.8000 1.0250 0.9000 1.4500 ;
    END
    ANTENNAGATEAREA 0.0582 ;
  END SE

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.4400 1.8000 1.5500 ;
    END
    ANTENNAGATEAREA 0.0666 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5550 1.3400 0.6450 ;
      RECT 1.2500 0.6450 1.3400 1.3550 ;
      RECT 0.0450 0.8150 0.7250 0.9050 ;
      RECT 0.6350 0.6450 0.7250 0.8150 ;
      RECT 0.0450 1.6950 0.1950 1.8800 ;
      RECT 0.0450 0.9050 0.1350 1.6950 ;
      RECT 1.2800 1.8300 1.9900 1.9200 ;
      RECT 2.1000 1.8750 2.2700 1.9650 ;
      RECT 2.1000 1.7400 2.1900 1.8750 ;
      RECT 0.8300 1.6500 2.1900 1.7400 ;
      RECT 2.0000 0.9100 2.0900 1.6500 ;
      RECT 1.8750 0.8200 2.0900 0.9100 ;
      RECT 1.8750 0.4800 1.9750 0.8200 ;
      RECT 0.8300 1.7400 0.9300 1.8800 ;
      RECT 0.9900 0.9100 1.0800 1.6500 ;
      RECT 0.8550 0.8100 1.0800 0.9100 ;
      RECT 2.3600 1.1300 3.1400 1.2300 ;
      RECT 2.3600 1.8700 2.5300 1.9700 ;
      RECT 2.3600 1.2300 2.4500 1.8700 ;
      RECT 2.3600 0.7450 2.4500 1.1300 ;
      RECT 2.8000 1.5350 3.3550 1.6250 ;
      RECT 2.8000 1.3250 2.8950 1.5350 ;
      RECT 3.2500 0.7050 3.3550 1.5350 ;
      RECT 3.4450 1.6250 4.2800 1.7150 ;
      RECT 4.1900 1.0100 4.2800 1.6250 ;
      RECT 3.4450 0.9300 3.5350 1.6250 ;
      RECT 3.4450 0.7450 3.6050 0.9300 ;
      RECT 4.3700 1.5500 4.5300 1.7400 ;
      RECT 4.4400 0.8900 4.5300 1.5500 ;
      RECT 3.8950 0.8000 4.5300 0.8900 ;
      RECT 3.8950 0.8900 3.9850 1.5300 ;
      RECT 5.0300 1.6500 5.2350 1.7400 ;
      RECT 5.0300 0.5950 5.1200 1.6500 ;
      RECT 5.0300 0.5700 5.2300 0.5950 ;
      RECT 2.1800 0.4800 5.2300 0.5700 ;
      RECT 2.1800 0.5700 2.2700 1.5400 ;
      RECT 3.6950 0.5700 3.7850 1.3600 ;
      RECT 3.4000 0.4200 3.5700 0.4800 ;
      RECT 3.6400 1.3600 3.7850 1.5300 ;
      RECT 3.1950 1.8300 5.7250 1.9200 ;
      RECT 5.3450 1.8200 5.7250 1.8300 ;
      RECT 5.6250 1.6500 5.7250 1.8200 ;
      RECT 5.2400 0.8200 5.7250 0.9100 ;
      RECT 5.6250 0.4150 5.7250 0.8200 ;
      RECT 5.3450 1.5400 5.4350 1.8200 ;
      RECT 5.2400 1.4500 5.4350 1.5400 ;
      RECT 5.2400 0.9100 5.3300 1.4500 ;
      RECT 3.3400 1.9200 3.5100 1.9900 ;
      RECT 3.1950 1.8150 3.2850 1.8300 ;
      RECT 2.6050 1.7250 3.2850 1.8150 ;
      RECT 2.6050 1.6100 2.6950 1.7250 ;
  END
END A2SDFFQN_X1M_A12TH

MACRO A2SDFFQN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6750 ;
        RECT 2.6800 0.3200 2.8900 0.3900 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9800 5.7500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.9750 0.5700 1.4200 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 3.8800 2.0100 4.0500 2.0800 ;
        RECT 2.7500 1.9000 2.8750 2.0800 ;
        RECT 0.3300 1.6850 0.4400 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 1.2000 1.9300 1.3050 ;
        RECT 1.6500 1.3050 1.7600 1.4850 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.1400 0.3500 1.5900 ;
    END
    ANTENNAGATEAREA 0.0654 ;
  END SE

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4100 1.0600 1.5500 1.4300 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END B

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 0.7800 4.9500 1.2900 ;
        RECT 4.7450 1.2900 4.9500 1.3900 ;
        RECT 4.6900 0.6800 4.9500 0.7800 ;
        RECT 4.7450 1.3900 4.8450 1.7200 ;
    END
    ANTENNADIFFAREA 0.323 ;
  END QN
  OBS
    LAYER M1 ;
      RECT 0.0500 0.7750 0.7800 0.8650 ;
      RECT 0.6900 0.8650 0.7800 1.4450 ;
      RECT 0.0500 1.7000 0.2000 1.8950 ;
      RECT 0.0500 0.8650 0.1400 1.7000 ;
      RECT 0.0500 0.5050 0.1800 0.7750 ;
      RECT 1.7050 1.9200 1.9050 1.9900 ;
      RECT 1.2000 1.9000 1.9050 1.9200 ;
      RECT 1.2000 1.8300 1.7950 1.9000 ;
      RECT 0.7850 1.6500 2.1100 1.7400 ;
      RECT 0.7600 0.5400 1.9750 0.6300 ;
      RECT 1.8850 0.6300 1.9750 0.9200 ;
      RECT 0.7850 1.7400 0.8850 1.8700 ;
      RECT 0.9350 0.6400 1.0250 1.6500 ;
      RECT 0.7600 0.6300 1.0250 0.6400 ;
      RECT 2.2450 1.1550 2.9300 1.2550 ;
      RECT 2.2200 1.7850 2.3350 1.9550 ;
      RECT 2.2450 1.2550 2.3350 1.7850 ;
      RECT 2.2450 0.7650 2.3350 1.1550 ;
      RECT 2.5500 1.4300 3.2400 1.5300 ;
      RECT 3.0300 0.6600 3.1300 1.3250 ;
      RECT 3.1450 1.5300 3.2400 1.7200 ;
      RECT 3.0300 1.3250 3.2400 1.5300 ;
      RECT 3.3400 1.6500 4.0500 1.7400 ;
      RECT 3.9600 1.1700 4.0500 1.6500 ;
      RECT 3.3400 0.6800 3.4350 1.6500 ;
      RECT 3.9600 1.0700 4.3600 1.1700 ;
      RECT 4.2300 1.6500 4.5600 1.7400 ;
      RECT 4.4700 0.8250 4.5600 1.6500 ;
      RECT 3.7700 0.7350 4.5600 0.8250 ;
      RECT 3.7700 0.8250 3.8600 1.1800 ;
      RECT 5.2150 1.5850 5.4300 1.6850 ;
      RECT 5.2150 0.5700 5.3050 1.5850 ;
      RECT 2.0650 0.4800 5.3050 0.5700 ;
      RECT 2.0650 0.5700 2.1550 1.4200 ;
      RECT 3.5500 0.5700 3.6400 1.4350 ;
      RECT 3.1800 0.4100 3.3500 0.4800 ;
      RECT 1.9800 1.4200 2.1550 1.5200 ;
      RECT 3.5500 1.4350 3.7450 1.5350 ;
      RECT 2.9650 1.8300 5.7700 1.9200 ;
      RECT 5.6800 1.6800 5.7700 1.8300 ;
      RECT 5.6800 1.5900 5.9550 1.6800 ;
      RECT 5.8650 0.5900 5.9550 1.5900 ;
      RECT 5.4000 0.5000 5.9550 0.5900 ;
      RECT 5.4000 0.5900 5.4900 1.1400 ;
      RECT 3.2350 1.9200 3.4050 1.9900 ;
      RECT 2.9650 1.7600 3.0550 1.8300 ;
      RECT 2.4350 1.6700 3.0550 1.7600 ;
      RECT 2.4350 1.7600 2.5250 1.8550 ;
  END
END A2SDFFQN_X2M_A12TH

MACRO A2SDFFQN_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4300 ;
        RECT 0.9850 0.3200 1.0850 0.6050 ;
        RECT 3.8150 0.3200 4.1850 0.3950 ;
        RECT 5.6950 0.3200 5.8150 0.6000 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.2150 0.9500 1.3900 ;
        RECT 0.7700 1.0150 0.9500 1.2150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.8800 5.1500 1.2500 ;
        RECT 4.6200 1.2500 5.2400 1.3500 ;
        RECT 4.5850 0.7800 5.2800 0.8800 ;
        RECT 4.6200 1.3500 4.7200 1.7250 ;
        RECT 5.1400 1.3500 5.2400 1.7250 ;
    END
    ANTENNADIFFAREA 0.5616 ;
  END QN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 1.0200 5.9500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 1.0600 1.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.0864 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0600 1.4250 1.3900 ;
    END
    ANTENNAGATEAREA 0.0864 ;
  END B

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0150 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 3.8150 2.0000 4.1850 2.0800 ;
        RECT 0.8700 1.7900 0.9800 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4850 0.4200 0.8000 0.5200 ;
      RECT 0.5800 1.9200 0.7500 1.9550 ;
      RECT 0.0500 1.8200 0.7500 1.9200 ;
      RECT 0.0500 0.5200 0.5850 0.6200 ;
      RECT 0.0500 0.6200 0.1500 1.8200 ;
      RECT 1.5650 1.9100 1.8450 1.9900 ;
      RECT 1.1150 1.9000 1.8450 1.9100 ;
      RECT 1.1150 1.8200 1.6550 1.9000 ;
      RECT 1.9000 1.6800 1.9900 1.7750 ;
      RECT 0.4400 1.5900 1.9900 1.6800 ;
      RECT 0.3700 0.8150 1.8700 0.9150 ;
      RECT 1.7700 0.4650 1.8700 0.8150 ;
      RECT 0.4400 0.9150 0.5300 1.5900 ;
      RECT 2.1000 1.6350 2.3200 1.7250 ;
      RECT 2.2300 0.9900 2.3200 1.6350 ;
      RECT 2.1550 0.8800 2.3200 0.9900 ;
      RECT 2.1550 0.7900 2.8650 0.8800 ;
      RECT 2.7750 0.8800 2.8650 1.2400 ;
      RECT 2.5300 1.6150 3.0600 1.7050 ;
      RECT 2.5300 1.0850 2.6200 1.6150 ;
      RECT 2.9700 0.7300 3.0600 1.6150 ;
      RECT 3.1500 1.4850 3.3800 1.5850 ;
      RECT 3.1500 0.9150 3.2500 1.4850 ;
      RECT 3.1500 0.8150 4.0050 0.9150 ;
      RECT 3.9050 0.9150 4.0050 1.0850 ;
      RECT 3.9050 1.0850 4.3150 1.1850 ;
      RECT 3.6650 1.4900 4.4950 1.5800 ;
      RECT 3.6650 1.0250 3.7550 1.4900 ;
      RECT 4.4050 0.9700 4.4950 1.4900 ;
      RECT 4.1800 0.8800 4.4950 0.9700 ;
      RECT 4.1800 0.8000 4.2700 0.8800 ;
      RECT 1.9750 0.4850 5.4850 0.5750 ;
      RECT 5.3950 0.5750 5.4850 1.7300 ;
      RECT 1.8800 1.4000 2.0650 1.5000 ;
      RECT 1.9750 0.5750 2.0650 1.4000 ;
      RECT 3.3500 0.4100 3.5200 0.4850 ;
      RECT 2.2800 1.8200 6.1550 1.9100 ;
      RECT 6.0650 0.7900 6.1550 1.8200 ;
      RECT 5.5900 0.7000 6.1550 0.7900 ;
      RECT 5.5900 0.7900 5.6800 1.2400 ;
      RECT 2.2800 1.9100 2.3900 1.9900 ;
      RECT 3.4350 1.9100 3.6350 1.9900 ;
      RECT 3.4700 1.1350 3.5600 1.8200 ;
      RECT 3.3450 1.0350 3.5600 1.1350 ;
  END
END A2SDFFQN_X3M_A12TH

MACRO A2SDFFQ_X0P5M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.6450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7400 ;
        RECT 1.0250 0.3200 1.1950 0.4350 ;
        RECT 2.6750 0.3200 2.8450 0.3900 ;
        RECT 3.8150 0.3200 3.9150 0.6750 ;
        RECT 5.1100 0.3200 5.2100 0.5750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8500 1.4100 5.0400 1.5900 ;
        RECT 4.9400 1.1600 5.0400 1.4100 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4500 0.7800 4.5500 1.2650 ;
        RECT 4.3550 1.2650 4.5500 1.3650 ;
        RECT 4.3800 0.6800 4.5500 0.7800 ;
        RECT 4.3550 1.3650 4.4750 1.7250 ;
    END
    ANTENNADIFFAREA 0.1668 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.3100 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.6450 2.7200 ;
        RECT 0.3300 1.8400 0.4400 2.0800 ;
        RECT 1.0550 1.8400 1.1650 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6500 0.7900 1.8250 1.1600 ;
    END
    ANTENNAGATEAREA 0.033 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2600 1.4500 0.9000 1.5500 ;
        RECT 0.2600 1.5500 0.3700 1.6650 ;
        RECT 0.8000 1.0050 0.9000 1.4500 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SE

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2100 1.4250 1.5200 1.5550 ;
        RECT 1.4300 1.1850 1.5200 1.4250 ;
    END
    ANTENNAGATEAREA 0.033 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5700 1.2600 0.6600 ;
      RECT 1.1700 0.6600 1.2600 0.8950 ;
      RECT 0.0700 0.8300 0.7250 0.9200 ;
      RECT 0.6350 0.6600 0.7250 0.8300 ;
      RECT 0.0700 1.8150 0.2100 1.9850 ;
      RECT 0.0700 0.9200 0.1600 1.8150 ;
      RECT 0.0700 0.6850 0.1800 0.8300 ;
      RECT 1.2750 1.8300 2.0250 1.9200 ;
      RECT 0.8350 1.6500 1.9750 1.7400 ;
      RECT 1.8850 1.6100 1.9750 1.6500 ;
      RECT 1.8850 1.5200 2.0750 1.6100 ;
      RECT 1.3700 0.5200 1.9350 0.6100 ;
      RECT 1.8350 0.4200 1.9350 0.5200 ;
      RECT 0.9900 1.0050 1.4600 1.0950 ;
      RECT 1.3700 0.6100 1.4600 1.0050 ;
      RECT 0.9900 1.0950 1.0800 1.6500 ;
      RECT 0.9900 0.8500 1.0800 1.0050 ;
      RECT 0.8800 0.7500 1.0800 0.8500 ;
      RECT 0.8350 1.7400 0.9250 1.9900 ;
      RECT 2.2250 1.2400 2.3150 1.7500 ;
      RECT 2.2250 1.1400 2.9600 1.2400 ;
      RECT 2.8600 1.2400 2.9600 1.3550 ;
      RECT 2.2250 0.6800 2.3150 1.1400 ;
      RECT 3.0500 1.5950 3.2200 1.6950 ;
      RECT 3.0500 1.0500 3.1400 1.5950 ;
      RECT 2.5450 0.9600 3.1400 1.0500 ;
      RECT 3.0300 0.8150 3.1400 0.9600 ;
      RECT 3.0300 0.7150 3.2250 0.8150 ;
      RECT 3.3200 1.6050 4.0200 1.7050 ;
      RECT 3.9200 1.1850 4.0200 1.6050 ;
      RECT 3.3200 0.6800 3.4200 1.6050 ;
      RECT 4.1300 1.0750 4.3600 1.1550 ;
      RECT 3.6950 0.9850 4.3600 1.0750 ;
      RECT 4.1300 1.1550 4.2300 1.7400 ;
      RECT 3.6950 1.0750 3.7850 1.1800 ;
      RECT 4.1850 0.6800 4.2850 0.9850 ;
      RECT 2.4200 1.8300 5.3400 1.9200 ;
      RECT 5.2500 0.9750 5.3400 1.8300 ;
      RECT 4.7500 0.8850 5.3400 0.9750 ;
      RECT 4.7500 0.6800 4.8400 0.8850 ;
      RECT 2.4200 1.3500 2.5100 1.8300 ;
      RECT 4.9300 0.6850 5.5200 0.7750 ;
      RECT 5.4300 0.7750 5.5200 1.9650 ;
      RECT 1.9450 1.2900 2.1350 1.3800 ;
      RECT 2.0450 0.5700 2.1350 1.2900 ;
      RECT 2.0450 0.4800 3.6050 0.5700 ;
      RECT 3.5150 0.5700 3.6050 0.7850 ;
      RECT 3.5150 0.8750 3.6050 1.4900 ;
      RECT 4.0050 0.4800 5.0200 0.5700 ;
      RECT 4.9300 0.5700 5.0200 0.6850 ;
      RECT 3.5150 0.7850 4.0950 0.8750 ;
      RECT 4.0050 0.5700 4.0950 0.7850 ;
  END
END A2SDFFQ_X0P5M_A12TH

MACRO A2SDFFQ_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.3550 0.3200 0.5250 0.7250 ;
        RECT 0.8850 0.3200 1.2550 0.3450 ;
        RECT 5.3400 0.3200 5.4500 0.6400 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4500 1.0100 5.6350 1.1900 ;
        RECT 5.5300 1.1900 5.6350 1.4150 ;
    END
    ANTENNAGATEAREA 0.0267 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6200 0.7250 4.7500 1.7100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4500 1.0100 0.6250 1.2000 ;
        RECT 0.4500 1.2000 0.5500 1.3500 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 0.8400 2.0600 1.2100 2.0800 ;
        RECT 3.8650 2.0200 4.2350 2.0800 ;
        RECT 2.9150 1.9050 3.0850 2.0800 ;
        RECT 0.3350 1.6900 0.4450 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4850 1.0500 1.9050 1.1500 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2500 1.4500 0.9000 1.5500 ;
        RECT 0.8000 1.0250 0.9000 1.4500 ;
    END
    ANTENNAGATEAREA 0.0618 ;
  END SE

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3900 1.4400 1.8500 1.5500 ;
    END
    ANTENNAGATEAREA 0.0726 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.6350 0.5550 1.3400 0.6450 ;
      RECT 1.2500 0.6450 1.3400 1.3550 ;
      RECT 0.0450 0.8150 0.7250 0.9050 ;
      RECT 0.6350 0.6450 0.7250 0.8150 ;
      RECT 0.0450 1.6950 0.1950 1.8800 ;
      RECT 0.0450 0.9050 0.1350 1.6950 ;
      RECT 1.2800 1.8300 1.9900 1.9200 ;
      RECT 2.1000 1.8750 2.2700 1.9650 ;
      RECT 2.1000 1.7400 2.1900 1.8750 ;
      RECT 0.8300 1.6500 2.1900 1.7400 ;
      RECT 2.0000 0.9100 2.0900 1.6500 ;
      RECT 1.8750 0.8200 2.0900 0.9100 ;
      RECT 1.8750 0.4800 1.9750 0.8200 ;
      RECT 0.8300 1.7400 0.9300 1.8800 ;
      RECT 0.9900 0.9100 1.0800 1.6500 ;
      RECT 0.8550 0.8100 1.0800 0.9100 ;
      RECT 2.3600 1.1300 3.1400 1.2300 ;
      RECT 2.3600 1.8700 2.5300 1.9700 ;
      RECT 2.3600 1.2300 2.4500 1.8700 ;
      RECT 2.3600 0.7450 2.4500 1.1300 ;
      RECT 2.8000 1.5200 3.3550 1.6150 ;
      RECT 2.8000 1.3250 2.8950 1.5200 ;
      RECT 3.2500 0.7200 3.3550 1.5200 ;
      RECT 3.4450 1.6250 4.2800 1.7150 ;
      RECT 4.1900 1.0900 4.2800 1.6250 ;
      RECT 3.4450 0.9300 3.5350 1.6250 ;
      RECT 3.4450 0.7450 3.6050 0.9300 ;
      RECT 4.3700 1.5500 4.5300 1.7400 ;
      RECT 4.4400 0.8450 4.5300 1.5500 ;
      RECT 3.8950 0.7550 4.5300 0.8450 ;
      RECT 3.8950 0.8450 3.9850 1.4050 ;
      RECT 5.0400 1.6500 5.2350 1.7400 ;
      RECT 5.0400 0.5950 5.1300 1.6500 ;
      RECT 5.0400 0.5700 5.2300 0.5950 ;
      RECT 2.1800 0.4800 5.2300 0.5700 ;
      RECT 2.1800 0.5700 2.2700 1.5400 ;
      RECT 3.6950 0.5700 3.7850 1.3600 ;
      RECT 3.4000 0.4200 3.5700 0.4800 ;
      RECT 3.6400 1.3600 3.7850 1.5300 ;
      RECT 3.1950 1.8300 5.7250 1.9200 ;
      RECT 5.3450 1.8200 5.7250 1.8300 ;
      RECT 5.6250 1.6500 5.7250 1.8200 ;
      RECT 5.2400 0.8200 5.7250 0.9100 ;
      RECT 5.6250 0.4150 5.7250 0.8200 ;
      RECT 5.3450 1.5400 5.4350 1.8200 ;
      RECT 5.2400 1.4500 5.4350 1.5400 ;
      RECT 5.2400 0.9100 5.3300 1.4500 ;
      RECT 3.3400 1.9200 3.5100 1.9900 ;
      RECT 3.1950 1.8150 3.2850 1.8300 ;
      RECT 2.6050 1.7250 3.2850 1.8150 ;
      RECT 2.6050 1.6100 2.6950 1.7250 ;
  END
END A2SDFFQ_X1M_A12TH

MACRO A2SDFFQ_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.0450 0.3200 ;
        RECT 0.3350 0.3200 0.4350 0.6750 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9800 5.7500 1.4100 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5000 1.2500 5.1250 1.3500 ;
        RECT 4.5000 1.3500 4.6000 1.7150 ;
        RECT 5.0250 1.3500 5.1250 1.7050 ;
        RECT 5.0250 0.7800 5.1250 1.2500 ;
        RECT 4.4000 0.6800 5.1250 0.7800 ;
    END
    ANTENNADIFFAREA 0.5088 ;
  END Q

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4450 0.9750 0.5700 1.4200 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.0450 2.7200 ;
        RECT 0.9250 2.0550 1.0950 2.0800 ;
        RECT 2.7750 2.0300 2.9900 2.0800 ;
        RECT 0.3300 1.6850 0.4400 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6100 1.2000 1.9300 1.3500 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.1400 0.3500 1.5900 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END SE

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0100 1.5250 1.1600 ;
        RECT 1.2500 1.1600 1.3500 1.2850 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END B
  OBS
    LAYER M1 ;
      RECT 0.0500 0.7750 0.7800 0.8650 ;
      RECT 0.6900 0.8650 0.7800 1.4450 ;
      RECT 0.0500 1.7000 0.2000 1.8950 ;
      RECT 0.0500 0.8650 0.1400 1.7000 ;
      RECT 0.0500 0.5050 0.1800 0.7750 ;
      RECT 1.7200 1.9200 1.8900 1.9650 ;
      RECT 1.2000 1.8300 1.8900 1.9200 ;
      RECT 0.7550 1.6500 2.1150 1.7400 ;
      RECT 0.9350 0.8100 1.9850 0.9000 ;
      RECT 1.8950 0.4800 1.9850 0.8100 ;
      RECT 0.7550 1.7400 0.9250 1.8150 ;
      RECT 0.9350 0.9000 1.0250 1.6500 ;
      RECT 0.9350 0.6400 1.0250 0.8100 ;
      RECT 0.7600 0.5400 1.0250 0.6400 ;
      RECT 2.2200 1.7600 2.3450 1.9700 ;
      RECT 2.2550 1.2550 2.3450 1.7600 ;
      RECT 2.2550 1.1550 2.9300 1.2550 ;
      RECT 2.2550 0.7650 2.3450 1.1550 ;
      RECT 3.1200 1.5250 3.2300 1.7400 ;
      RECT 2.5500 1.4250 3.2300 1.5250 ;
      RECT 3.0300 1.3700 3.2300 1.4250 ;
      RECT 3.0300 0.6600 3.1300 1.3700 ;
      RECT 3.3400 1.6500 4.1100 1.7400 ;
      RECT 4.0200 0.9700 4.1100 1.6500 ;
      RECT 3.3400 0.6800 3.4350 1.6500 ;
      RECT 4.2000 1.0400 4.9350 1.1400 ;
      RECT 4.2550 1.1400 4.3450 1.7200 ;
      RECT 4.2000 0.7700 4.2900 1.0400 ;
      RECT 3.7900 0.6800 4.2900 0.7700 ;
      RECT 3.7900 0.7700 3.8800 1.1800 ;
      RECT 5.2200 1.5850 5.4300 1.6850 ;
      RECT 5.2200 0.5700 5.3100 1.5850 ;
      RECT 2.0750 0.4800 5.3100 0.5700 ;
      RECT 2.0750 0.5700 2.1650 1.4200 ;
      RECT 3.5500 0.5700 3.6400 1.4350 ;
      RECT 3.1800 0.4100 3.3500 0.4800 ;
      RECT 1.9900 1.4200 2.1650 1.5200 ;
      RECT 3.5500 1.4350 3.7650 1.5350 ;
      RECT 2.4350 1.8300 5.7700 1.9200 ;
      RECT 5.6800 1.6800 5.7700 1.8300 ;
      RECT 5.6800 1.5900 5.9550 1.6800 ;
      RECT 5.8650 0.5900 5.9550 1.5900 ;
      RECT 5.4000 0.5000 5.9550 0.5900 ;
      RECT 5.4000 0.5900 5.4900 1.1400 ;
      RECT 3.2350 1.9200 3.4050 1.9900 ;
      RECT 2.4350 1.6700 2.5250 1.8300 ;
  END
END A2SDFFQ_X2M_A12TH

MACRO A2SDFFQ_X3M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4300 ;
        RECT 0.9850 0.3200 1.0850 0.6050 ;
        RECT 3.7350 0.3200 3.9050 0.3450 ;
        RECT 4.3050 0.3200 4.5200 0.3600 ;
        RECT 4.8200 0.3200 5.0350 0.3600 ;
        RECT 5.6950 0.3200 5.8150 0.6000 ;
    END
  END VSS

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8500 1.0200 5.9500 1.5000 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END CK

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8500 1.1950 0.9500 1.3900 ;
        RECT 0.7700 1.0150 0.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0500 0.9000 5.1500 1.2900 ;
        RECT 4.6200 1.2900 5.2400 1.3900 ;
        RECT 4.5650 0.8000 5.2850 0.9000 ;
        RECT 4.6200 1.3900 4.7200 1.7000 ;
        RECT 5.1400 1.3900 5.2400 1.7000 ;
    END
    ANTENNADIFFAREA 0.6048 ;
  END Q

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6000 1.0600 1.7500 1.3900 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2500 1.0600 1.4250 1.3900 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END B

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0150 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0678 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 0.8900 1.8300 0.9900 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.4000 0.4200 0.7800 0.5200 ;
      RECT 0.0500 1.8200 0.7650 1.9200 ;
      RECT 0.0500 0.5700 0.5000 0.6700 ;
      RECT 0.4000 0.5200 0.5000 0.5700 ;
      RECT 0.0500 0.6700 0.1500 1.8200 ;
      RECT 1.6900 1.9100 1.7900 1.9900 ;
      RECT 1.1150 1.8200 1.7900 1.9100 ;
      RECT 1.8950 1.6800 1.9850 1.7700 ;
      RECT 0.4400 1.5900 1.9850 1.6800 ;
      RECT 0.3700 0.8100 1.8700 0.9100 ;
      RECT 1.7700 0.4650 1.8700 0.8100 ;
      RECT 0.4400 0.9100 0.5300 1.5900 ;
      RECT 2.0950 1.6350 2.3150 1.7250 ;
      RECT 2.2250 0.9800 2.3150 1.6350 ;
      RECT 2.1400 0.8800 2.3150 0.9800 ;
      RECT 2.1400 0.7900 2.8600 0.8800 ;
      RECT 2.7700 0.8800 2.8600 1.2400 ;
      RECT 2.5250 1.6150 3.0550 1.7050 ;
      RECT 2.5250 1.0850 2.6150 1.6150 ;
      RECT 2.9650 0.7300 3.0550 1.6150 ;
      RECT 3.1700 1.4850 3.3800 1.5850 ;
      RECT 3.1700 0.9250 3.2700 1.4850 ;
      RECT 3.1700 0.8250 4.0050 0.9250 ;
      RECT 3.9050 0.9250 4.0050 1.2300 ;
      RECT 4.0950 1.0800 4.9550 1.1800 ;
      RECT 4.0950 1.4450 4.1950 1.7050 ;
      RECT 3.6750 1.3450 4.1950 1.4450 ;
      RECT 4.0950 1.1800 4.1950 1.3450 ;
      RECT 3.6750 1.0350 3.7750 1.3450 ;
      RECT 4.0950 0.7650 4.1950 1.0800 ;
      RECT 1.9600 0.4850 5.4850 0.5750 ;
      RECT 5.3950 0.5750 5.4850 1.7300 ;
      RECT 1.8650 1.3950 2.0500 1.4950 ;
      RECT 1.9600 0.5750 2.0500 1.3950 ;
      RECT 3.3500 0.4100 3.5200 0.4850 ;
      RECT 2.2750 1.8200 6.1550 1.9100 ;
      RECT 6.0650 0.7900 6.1550 1.8200 ;
      RECT 5.5900 0.7000 6.1550 0.7900 ;
      RECT 5.5900 0.7900 5.6800 1.2400 ;
      RECT 2.2750 1.9100 2.3850 1.9900 ;
      RECT 3.4350 1.9100 3.6350 1.9900 ;
      RECT 3.4700 1.1350 3.5600 1.8200 ;
      RECT 3.3600 1.0350 3.5600 1.1350 ;
  END
END A2SDFFQ_X3M_A12TH

MACRO A2SDFFQ_X4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.6450 0.3200 ;
        RECT 0.0450 0.3200 0.2150 0.4300 ;
        RECT 1.0000 0.3200 1.1000 0.5800 ;
        RECT 3.8150 0.3200 3.9850 0.3450 ;
        RECT 6.0900 0.3200 6.2000 0.7150 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7500 1.4400 5.4150 1.5600 ;
        RECT 4.7500 1.5600 4.8700 1.6650 ;
        RECT 5.2850 1.5600 5.4150 1.6800 ;
        RECT 4.7500 1.2900 4.8700 1.4400 ;
        RECT 5.2850 0.8900 5.4150 1.4400 ;
        RECT 4.7250 0.7700 5.4150 0.8900 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END Q

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1000 1.2400 1.5000 1.3550 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END B

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8300 1.0350 0.9500 1.4000 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2450 1.0200 6.3650 1.5000 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END CK

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3700 1.0500 1.7900 1.1500 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END A

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2400 1.0150 0.3500 1.4500 ;
    END
    ANTENNAGATEAREA 0.0696 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.6450 2.7200 ;
        RECT 0.8700 1.8400 0.9700 2.0800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 0.5750 1.9200 0.7450 1.9700 ;
      RECT 0.0500 1.8200 0.7450 1.9200 ;
      RECT 0.0500 0.5700 0.4950 0.6700 ;
      RECT 0.3950 0.5150 0.4950 0.5700 ;
      RECT 0.3950 0.4150 0.7750 0.5150 ;
      RECT 0.0500 0.6700 0.1500 1.8200 ;
      RECT 1.6900 1.9150 1.7900 1.9900 ;
      RECT 1.1150 1.8150 1.7900 1.9150 ;
      RECT 1.9450 1.6350 2.0350 1.9400 ;
      RECT 0.4600 1.5450 2.0350 1.6350 ;
      RECT 0.4600 0.7800 1.8700 0.8800 ;
      RECT 1.7700 0.4550 1.8700 0.7800 ;
      RECT 0.4600 0.8800 0.5500 1.5450 ;
      RECT 2.2000 0.8750 2.3000 1.6750 ;
      RECT 2.1550 0.7750 2.3000 0.8750 ;
      RECT 2.1550 0.6850 2.9750 0.7750 ;
      RECT 2.8850 0.7750 2.9750 1.2400 ;
      RECT 2.5400 1.5450 3.1550 1.6350 ;
      RECT 2.5400 1.0200 2.6300 1.5450 ;
      RECT 3.0650 0.7300 3.1550 1.5450 ;
      RECT 4.0200 1.2000 4.4550 1.3000 ;
      RECT 4.0200 0.9300 4.1200 1.2000 ;
      RECT 3.2550 0.8300 4.1200 0.9300 ;
      RECT 3.2550 0.9300 3.3550 1.7050 ;
      RECT 4.5450 1.0800 5.1850 1.1800 ;
      RECT 3.8300 1.5800 4.6350 1.6700 ;
      RECT 4.5450 1.1800 4.6350 1.5800 ;
      RECT 3.8300 1.0450 3.9200 1.5800 ;
      RECT 4.5450 0.9250 4.6350 1.0800 ;
      RECT 4.2300 0.8350 4.6350 0.9250 ;
      RECT 4.2300 0.7550 4.3200 0.8350 ;
      RECT 1.9600 0.4850 5.8850 0.5750 ;
      RECT 5.7950 0.5750 5.8850 1.7200 ;
      RECT 1.8800 1.3050 2.0500 1.4050 ;
      RECT 1.9600 0.5750 2.0500 1.3050 ;
      RECT 3.5150 0.4100 3.6850 0.4850 ;
      RECT 2.3450 1.8150 6.5550 1.9050 ;
      RECT 6.4650 0.9050 6.5550 1.8150 ;
      RECT 5.9800 0.8150 6.5550 0.9050 ;
      RECT 6.4250 0.5200 6.5550 0.8150 ;
      RECT 5.9800 0.9050 6.0700 1.4600 ;
      RECT 2.3450 1.9050 2.4650 1.9900 ;
      RECT 3.7650 1.9050 3.9100 1.9900 ;
      RECT 3.5950 1.0350 3.6950 1.8150 ;
  END
END A2SDFFQ_X4M_A12TH

MACRO ADDFCIN_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 4.7900 1.9250 4.9600 2.0800 ;
        RECT 5.3050 1.8300 5.4750 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 1.1900 1.1600 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.4000 0.3200 0.6100 0.3600 ;
        RECT 4.6750 0.3200 4.8550 0.3300 ;
    END
  END VSS

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9100 5.7500 1.4900 ;
        RECT 5.6000 1.4900 5.7500 1.5900 ;
        RECT 5.6000 0.8100 5.7500 0.9100 ;
        RECT 5.6000 1.5900 5.7000 1.9800 ;
        RECT 5.6000 0.4800 5.7000 0.8100 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END SUM

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7800 2.7500 1.2500 ;
        RECT 2.6500 1.2500 3.0400 1.3800 ;
        RECT 2.6500 0.6600 3.0400 0.7800 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END CO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.0650 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2352 ;
  END B

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6100 0.8100 4.7900 1.1950 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END CIN
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5550 0.5700 ;
      RECT 0.0450 1.4500 0.1750 1.8300 ;
      RECT 0.0450 0.8850 0.1350 1.4500 ;
      RECT 0.0450 0.5700 0.1750 0.8850 ;
      RECT 0.0450 1.8300 1.2750 1.9200 ;
      RECT 0.2650 0.6600 1.9800 0.7500 ;
      RECT 1.8900 0.7500 1.9800 1.3450 ;
      RECT 1.8800 0.6100 1.9800 0.6600 ;
      RECT 1.8550 1.3450 1.9800 1.5400 ;
      RECT 1.8800 0.5100 2.2400 0.6100 ;
      RECT 0.2650 1.6450 0.7350 1.7350 ;
      RECT 0.2650 1.2400 0.3550 1.6450 ;
      RECT 0.2350 0.9950 0.3550 1.2400 ;
      RECT 0.2650 0.7500 0.3550 0.9950 ;
      RECT 2.1000 1.4700 3.4300 1.5600 ;
      RECT 3.1850 1.4500 3.4300 1.4700 ;
      RECT 2.3800 0.4800 3.4200 0.5700 ;
      RECT 3.2450 0.4600 3.4200 0.4800 ;
      RECT 2.1000 0.8050 2.2000 1.4700 ;
      RECT 2.1000 0.7150 2.4700 0.8050 ;
      RECT 2.3800 0.5700 2.4700 0.7150 ;
      RECT 3.5400 1.3150 3.6500 1.4650 ;
      RECT 3.1300 1.2150 3.6500 1.3150 ;
      RECT 3.1300 1.0850 3.2200 1.2150 ;
      RECT 2.8450 0.9850 3.2200 1.0850 ;
      RECT 3.1300 0.7700 3.2200 0.9850 ;
      RECT 3.1300 0.6700 3.6400 0.7700 ;
      RECT 3.5350 0.4300 3.6400 0.6700 ;
      RECT 1.3050 1.4700 1.7450 1.5600 ;
      RECT 1.5900 0.8400 1.7950 0.9500 ;
      RECT 1.6550 1.5600 1.7450 1.6500 ;
      RECT 1.6550 0.9500 1.7450 1.4700 ;
      RECT 1.6550 1.6500 3.8700 1.7400 ;
      RECT 3.3150 0.8650 3.9900 0.9850 ;
      RECT 3.7700 1.1050 3.8700 1.6500 ;
      RECT 3.7700 0.8650 3.9900 1.1050 ;
      RECT 3.2950 1.9200 3.5100 1.9900 ;
      RECT 1.3950 1.9000 4.3100 1.9200 ;
      RECT 4.0100 1.9200 4.3100 1.9900 ;
      RECT 1.3950 1.8300 4.1150 1.9000 ;
      RECT 1.3950 1.7400 1.4850 1.8300 ;
      RECT 0.8550 1.6500 1.4850 1.7400 ;
      RECT 0.4550 0.9300 0.5450 1.4450 ;
      RECT 0.8550 1.5350 0.9450 1.6500 ;
      RECT 0.4550 1.4450 0.9450 1.5350 ;
      RECT 0.4550 0.8400 1.2800 0.9300 ;
      RECT 4.2700 1.2900 5.1500 1.3800 ;
      RECT 5.0600 1.0200 5.1500 1.2900 ;
      RECT 4.2700 0.7700 4.3700 1.2900 ;
      RECT 4.2700 0.6600 4.4700 0.7700 ;
      RECT 3.9950 1.4700 5.3300 1.5600 ;
      RECT 5.2400 0.7500 5.3300 1.4700 ;
      RECT 5.0250 0.6600 5.3300 0.7500 ;
      RECT 3.9950 1.5600 4.1150 1.6750 ;
      RECT 3.9950 1.2700 4.1800 1.4700 ;
      RECT 4.0800 0.7700 4.1800 1.2700 ;
      RECT 3.7950 0.6700 4.1800 0.7700 ;
      RECT 3.7950 0.4300 3.9050 0.6700 ;
      RECT 4.2450 1.6500 5.5100 1.7400 ;
      RECT 5.4200 0.5700 5.5100 1.6500 ;
      RECT 4.0250 0.4800 5.5100 0.5700 ;
      RECT 4.0250 0.4600 4.2500 0.4800 ;
  END
END ADDFCIN_X1M_A12TH

MACRO ADDFCIN_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.5800 2.0100 2.7900 2.0800 ;
        RECT 3.1200 2.0100 3.3300 2.0800 ;
        RECT 4.9350 1.9750 5.1050 2.0800 ;
        RECT 5.4700 1.9650 5.6000 2.0800 ;
        RECT 6.0050 1.7600 6.1050 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 1.1900 1.1600 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4000 0.3200 0.6100 0.3600 ;
        RECT 2.5800 0.3200 2.7900 0.3900 ;
        RECT 3.1200 0.3200 3.3100 0.3900 ;
        RECT 6.0050 0.3200 6.1050 0.6400 ;
    END
  END VSS

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7450 1.4500 6.1500 1.5500 ;
        RECT 5.7450 1.5500 5.8450 1.9800 ;
        RECT 6.0500 0.9500 6.1500 1.4500 ;
        RECT 5.7450 0.8500 6.1500 0.9500 ;
        RECT 5.7450 0.4800 5.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END SUM

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7600 2.7500 1.2500 ;
        RECT 2.6500 1.2500 3.0550 1.3800 ;
        RECT 2.6500 0.6600 3.0550 0.7600 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END CO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.0700 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2412 ;
  END B

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8050 0.8100 4.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0945 ;
  END CIN
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5550 0.5700 ;
      RECT 0.0450 1.4500 0.1750 1.8300 ;
      RECT 0.0450 0.8850 0.1350 1.4500 ;
      RECT 0.0450 0.5700 0.1750 0.8850 ;
      RECT 0.0450 1.8300 1.2750 1.9200 ;
      RECT 0.2650 0.6600 1.9800 0.7500 ;
      RECT 1.8900 0.7500 1.9800 1.3450 ;
      RECT 1.8800 0.6100 1.9800 0.6600 ;
      RECT 1.8550 1.3450 1.9800 1.5400 ;
      RECT 1.8800 0.5100 2.2400 0.6100 ;
      RECT 0.2650 1.6450 0.7450 1.7350 ;
      RECT 0.2650 1.2400 0.3550 1.6450 ;
      RECT 0.2350 0.9950 0.3550 1.2400 ;
      RECT 0.2650 0.7500 0.3550 0.9950 ;
      RECT 2.1000 1.4700 3.5750 1.5600 ;
      RECT 3.3300 1.4500 3.5750 1.4700 ;
      RECT 2.3800 0.4800 3.5650 0.5700 ;
      RECT 3.3900 0.4600 3.5650 0.4800 ;
      RECT 2.1000 0.8050 2.2000 1.4700 ;
      RECT 2.1000 0.7150 2.4700 0.8050 ;
      RECT 2.3800 0.5700 2.4700 0.7150 ;
      RECT 3.6850 1.3150 3.7850 1.5500 ;
      RECT 3.1900 1.2150 3.7850 1.3150 ;
      RECT 3.1900 1.0850 3.2900 1.2150 ;
      RECT 2.9050 0.9850 3.2900 1.0850 ;
      RECT 3.1900 0.7700 3.2900 0.9850 ;
      RECT 3.1900 0.6700 3.7900 0.7700 ;
      RECT 3.6800 0.4300 3.7900 0.6700 ;
      RECT 1.3050 1.4700 1.7450 1.5600 ;
      RECT 1.5900 0.8400 1.7950 0.9500 ;
      RECT 1.6550 1.5600 1.7450 1.6500 ;
      RECT 1.6550 0.9500 1.7450 1.4700 ;
      RECT 1.6550 1.6500 4.0150 1.7400 ;
      RECT 3.4600 0.8650 4.1350 0.9650 ;
      RECT 3.9150 1.1050 4.0150 1.6500 ;
      RECT 3.9150 0.8650 4.1350 1.1050 ;
      RECT 3.4450 1.9200 3.6550 1.9900 ;
      RECT 1.3950 1.9000 4.4550 1.9200 ;
      RECT 4.1650 1.9200 4.4550 1.9900 ;
      RECT 1.3950 1.8300 4.2700 1.9000 ;
      RECT 1.3950 1.7400 1.4850 1.8300 ;
      RECT 0.8550 1.6500 1.4850 1.7400 ;
      RECT 0.4550 0.9300 0.5450 1.4450 ;
      RECT 0.8550 1.5350 0.9450 1.6500 ;
      RECT 0.4550 1.4450 0.9450 1.5350 ;
      RECT 0.4550 0.8400 1.2800 0.9300 ;
      RECT 4.4150 1.3400 5.2250 1.4300 ;
      RECT 5.1350 0.9900 5.2250 1.3400 ;
      RECT 4.4150 0.7700 4.5150 1.3400 ;
      RECT 4.4150 0.6600 4.6150 0.7700 ;
      RECT 4.1400 1.5200 5.4750 1.6100 ;
      RECT 5.3850 0.7500 5.4750 1.5200 ;
      RECT 5.1700 0.6600 5.4750 0.7500 ;
      RECT 4.1400 1.6100 4.2600 1.6750 ;
      RECT 4.1400 1.2700 4.3250 1.5200 ;
      RECT 4.2250 0.7700 4.3250 1.2700 ;
      RECT 3.9400 0.6700 4.3250 0.7700 ;
      RECT 3.9400 0.4300 4.0450 0.6700 ;
      RECT 5.5650 1.0500 5.8550 1.1500 ;
      RECT 4.3900 1.7000 5.6550 1.7900 ;
      RECT 5.5650 1.1500 5.6550 1.7000 ;
      RECT 5.5650 0.5700 5.6550 1.0500 ;
      RECT 4.1700 0.4800 5.6550 0.5700 ;
      RECT 4.1700 0.4600 4.3950 0.4800 ;
  END
END ADDFCIN_X1P4M_A12TH

MACRO ADDFCIN_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.6200 2.0450 2.7900 2.0800 ;
        RECT 3.1400 2.0450 3.3100 2.0800 ;
        RECT 4.9350 2.0350 5.1050 2.0800 ;
        RECT 5.4500 1.8700 5.6200 2.0800 ;
        RECT 6.0050 1.7600 6.1050 2.0800 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 1.1900 1.1600 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4000 0.3200 0.6100 0.3600 ;
        RECT 6.0050 0.3200 6.1050 0.6400 ;
    END
  END VSS

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7450 1.2500 6.1500 1.3500 ;
        RECT 5.7450 1.3500 5.8450 1.7150 ;
        RECT 6.0500 0.9500 6.1500 1.2500 ;
        RECT 5.7450 0.8500 6.1500 0.9500 ;
        RECT 5.7450 0.4300 5.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END SUM

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7600 2.7500 1.2500 ;
        RECT 2.6500 1.2500 3.0800 1.3800 ;
        RECT 2.6500 0.6600 3.0800 0.7600 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END CO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.0750 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2451 ;
  END B

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8050 0.8100 4.9500 1.1950 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END CIN
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5550 0.5700 ;
      RECT 0.0450 1.4500 0.1750 1.8300 ;
      RECT 0.0450 0.8850 0.1350 1.4500 ;
      RECT 0.0450 0.5700 0.1750 0.8850 ;
      RECT 0.0450 1.8300 1.2750 1.9200 ;
      RECT 0.2650 0.6600 1.9800 0.7500 ;
      RECT 1.8900 0.7500 1.9800 1.3450 ;
      RECT 1.8800 0.6100 1.9800 0.6600 ;
      RECT 1.8550 1.3450 1.9800 1.5400 ;
      RECT 1.8800 0.5100 2.2400 0.6100 ;
      RECT 0.2650 1.6450 0.7350 1.7350 ;
      RECT 0.2650 1.2400 0.3550 1.6450 ;
      RECT 0.2350 0.9950 0.3550 1.2400 ;
      RECT 0.2650 0.7500 0.3550 0.9950 ;
      RECT 2.1000 1.4700 3.5750 1.5600 ;
      RECT 3.3300 1.4500 3.5750 1.4700 ;
      RECT 2.4000 0.4800 3.5650 0.5700 ;
      RECT 3.3400 0.4600 3.5650 0.4800 ;
      RECT 2.1000 0.8050 2.2000 1.4700 ;
      RECT 2.1000 0.7150 2.4900 0.8050 ;
      RECT 2.4000 0.5700 2.4900 0.7150 ;
      RECT 3.6850 1.3150 3.7850 1.5500 ;
      RECT 3.1900 1.2150 3.7850 1.3150 ;
      RECT 3.1900 1.0850 3.2900 1.2150 ;
      RECT 2.9050 0.9850 3.2900 1.0850 ;
      RECT 3.1900 0.7700 3.2900 0.9850 ;
      RECT 3.1900 0.6700 3.7900 0.7700 ;
      RECT 3.6800 0.4300 3.7900 0.6700 ;
      RECT 1.3050 1.4700 1.7450 1.5600 ;
      RECT 1.5900 0.8400 1.7950 0.9500 ;
      RECT 1.6550 1.5600 1.7450 1.6500 ;
      RECT 1.6550 0.9500 1.7450 1.4700 ;
      RECT 1.6550 1.6500 4.0150 1.7400 ;
      RECT 3.4250 0.8650 4.1350 0.9650 ;
      RECT 3.9150 1.1050 4.0150 1.6500 ;
      RECT 3.9150 0.8650 4.1350 1.1050 ;
      RECT 3.4400 1.9200 3.6550 1.9900 ;
      RECT 1.3950 1.9000 4.4400 1.9200 ;
      RECT 4.1550 1.9200 4.4400 1.9900 ;
      RECT 1.3950 1.8300 4.2600 1.9000 ;
      RECT 1.3950 1.7400 1.4850 1.8300 ;
      RECT 0.8550 1.6500 1.4850 1.7400 ;
      RECT 0.4550 0.9300 0.5450 1.4450 ;
      RECT 0.8550 1.5350 0.9450 1.6500 ;
      RECT 0.4550 1.4450 0.9450 1.5350 ;
      RECT 0.4550 0.8400 1.2800 0.9300 ;
      RECT 4.4150 1.3300 5.2250 1.4200 ;
      RECT 5.1350 0.9900 5.2250 1.3300 ;
      RECT 4.4150 0.7700 4.5150 1.3300 ;
      RECT 4.4150 0.6600 4.6150 0.7700 ;
      RECT 4.1400 1.5100 5.4750 1.6000 ;
      RECT 5.3850 0.7500 5.4750 1.5100 ;
      RECT 5.1700 0.6600 5.4750 0.7500 ;
      RECT 4.1400 1.6000 4.2600 1.6750 ;
      RECT 4.1400 1.2700 4.3250 1.5100 ;
      RECT 4.2250 0.7700 4.3250 1.2700 ;
      RECT 3.9400 0.6700 4.3250 0.7700 ;
      RECT 3.9400 0.4300 4.0500 0.6700 ;
      RECT 5.5650 1.0500 5.8550 1.1500 ;
      RECT 4.3700 1.6900 5.6550 1.7800 ;
      RECT 5.5650 1.1500 5.6550 1.6900 ;
      RECT 5.5650 0.5700 5.6550 1.0500 ;
      RECT 4.1700 0.4800 5.6550 0.5700 ;
      RECT 4.1700 0.4600 4.3950 0.4800 ;
  END
END ADDFCIN_X2M_A12TH

MACRO ADDFH_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 5.8450 2.7200 ;
        RECT 4.7900 1.9250 4.9600 2.0800 ;
        RECT 5.3050 1.8750 5.4750 2.0800 ;
    END
  END VDD

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.0100 0.8500 5.1900 1.2150 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END CI

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.0650 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2352 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 5.8450 0.3200 ;
        RECT 0.4000 0.3200 0.6100 0.3600 ;
        RECT 4.6750 0.3200 4.8550 0.3300 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7800 2.7500 1.2500 ;
        RECT 2.6500 1.2500 3.0400 1.3800 ;
        RECT 2.6500 0.6600 3.0400 0.7800 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END CO

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.6500 0.9100 5.7500 1.3100 ;
        RECT 5.6200 1.3100 5.7500 1.4100 ;
        RECT 5.6200 0.8100 5.7500 0.9100 ;
        RECT 5.6200 1.4100 5.7200 1.8000 ;
        RECT 5.6200 0.4800 5.7200 0.8100 ;
    END
    ANTENNADIFFAREA 0.2925 ;
  END SUM

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 1.1900 1.1600 ;
    END
    ANTENNAGATEAREA 0.0876 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5550 0.5700 ;
      RECT 0.0450 1.4500 0.1750 1.8300 ;
      RECT 0.0450 0.8850 0.1350 1.4500 ;
      RECT 0.0450 0.5700 0.1750 0.8850 ;
      RECT 0.0450 1.8300 1.2750 1.9200 ;
      RECT 0.2650 0.6600 1.9800 0.7500 ;
      RECT 1.8900 0.7500 1.9800 1.3450 ;
      RECT 1.8800 0.6100 1.9800 0.6600 ;
      RECT 1.8550 1.3450 1.9800 1.5400 ;
      RECT 1.8800 0.5100 2.2400 0.6100 ;
      RECT 0.2650 1.6450 0.7350 1.7350 ;
      RECT 0.2650 1.2400 0.3550 1.6450 ;
      RECT 0.2350 0.9950 0.3550 1.2400 ;
      RECT 0.2650 0.7500 0.3550 0.9950 ;
      RECT 2.1000 1.4700 3.4300 1.5600 ;
      RECT 3.1850 1.4500 3.4300 1.4700 ;
      RECT 2.3800 0.4800 3.4200 0.5700 ;
      RECT 3.2450 0.4600 3.4200 0.4800 ;
      RECT 2.1000 0.8050 2.2000 1.4700 ;
      RECT 2.1000 0.7150 2.4700 0.8050 ;
      RECT 2.3800 0.5700 2.4700 0.7150 ;
      RECT 3.5400 1.3150 3.6500 1.4650 ;
      RECT 3.1300 1.2150 3.6500 1.3150 ;
      RECT 3.1300 1.0850 3.2200 1.2150 ;
      RECT 2.8450 0.9850 3.2200 1.0850 ;
      RECT 3.1300 0.7700 3.2200 0.9850 ;
      RECT 3.1300 0.6700 3.6450 0.7700 ;
      RECT 3.5350 0.4300 3.6450 0.6700 ;
      RECT 1.3050 1.4700 1.7450 1.5600 ;
      RECT 1.5900 0.8400 1.7950 0.9500 ;
      RECT 1.6550 1.5600 1.7450 1.6500 ;
      RECT 1.6550 0.9500 1.7450 1.4700 ;
      RECT 1.6550 1.6500 3.8700 1.7400 ;
      RECT 3.3150 0.8650 3.9900 0.9850 ;
      RECT 3.7700 1.1050 3.8700 1.6500 ;
      RECT 3.7700 0.8650 3.9900 1.1050 ;
      RECT 3.2950 1.9200 3.5100 1.9900 ;
      RECT 1.3950 1.9000 4.2900 1.9200 ;
      RECT 4.0100 1.9200 4.2900 1.9900 ;
      RECT 1.3950 1.8300 4.1150 1.9000 ;
      RECT 1.3950 1.7400 1.4850 1.8300 ;
      RECT 0.8550 1.6500 1.4850 1.7400 ;
      RECT 0.4550 0.9300 0.5450 1.4450 ;
      RECT 0.8550 1.5350 0.9450 1.6500 ;
      RECT 0.4550 1.4450 0.9450 1.5350 ;
      RECT 0.4550 0.8400 1.2800 0.9300 ;
      RECT 4.2750 1.3150 4.7200 1.4250 ;
      RECT 4.2750 0.7700 4.3750 1.3150 ;
      RECT 4.2750 0.6600 4.4850 0.7700 ;
      RECT 3.9950 1.5150 5.2400 1.6050 ;
      RECT 4.6700 0.6600 5.2250 0.7500 ;
      RECT 3.9950 1.6050 4.1150 1.6750 ;
      RECT 3.9950 1.2700 4.1800 1.5150 ;
      RECT 4.8250 1.1950 4.9150 1.5150 ;
      RECT 4.0800 0.7700 4.1800 1.2700 ;
      RECT 4.6700 1.1050 4.9150 1.1950 ;
      RECT 3.7950 0.6700 4.1800 0.7700 ;
      RECT 4.6700 0.7500 4.7600 1.1050 ;
      RECT 3.7950 0.4300 3.9050 0.6700 ;
      RECT 4.2450 1.6950 5.5300 1.7850 ;
      RECT 5.4400 0.5700 5.5300 1.6950 ;
      RECT 4.0250 0.4800 5.5300 0.5700 ;
      RECT 4.0250 0.4600 4.2500 0.4800 ;
  END
END ADDFH_X1M_A12TH

MACRO ADDFH_X1P4M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.5800 2.0100 2.7900 2.0800 ;
        RECT 3.1200 2.0100 3.3300 2.0800 ;
        RECT 4.9350 1.9750 5.1050 2.0800 ;
        RECT 5.4700 1.9650 5.6000 2.0800 ;
        RECT 6.0050 1.7600 6.1050 2.0800 ;
    END
  END VDD

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2350 0.9800 5.3900 1.2100 ;
        RECT 5.0100 0.8500 5.3900 0.9800 ;
    END
    ANTENNAGATEAREA 0.0945 ;
  END CI

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.0700 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2412 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4000 0.3200 0.6100 0.3600 ;
        RECT 2.5800 0.3200 2.7900 0.3900 ;
        RECT 3.1200 0.3200 3.3100 0.3900 ;
        RECT 6.0050 0.3200 6.1050 0.6400 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7600 2.7500 1.2500 ;
        RECT 2.6500 1.2500 3.0550 1.3800 ;
        RECT 2.6500 0.6600 3.0550 0.7600 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END CO

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7450 1.4500 6.1500 1.5500 ;
        RECT 5.7450 1.5500 5.8450 1.9800 ;
        RECT 6.0500 0.9500 6.1500 1.4500 ;
        RECT 5.7450 0.8500 6.1500 0.9500 ;
        RECT 5.7450 0.4800 5.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.231 ;
  END SUM

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 1.1900 1.1600 ;
    END
    ANTENNAGATEAREA 0.0936 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5550 0.5700 ;
      RECT 0.0450 1.4500 0.1750 1.8300 ;
      RECT 0.0450 0.8850 0.1350 1.4500 ;
      RECT 0.0450 0.5700 0.1750 0.8850 ;
      RECT 0.0450 1.8300 1.2750 1.9200 ;
      RECT 0.2650 0.6600 1.9800 0.7500 ;
      RECT 1.8900 0.7500 1.9800 1.3450 ;
      RECT 1.8800 0.6100 1.9800 0.6600 ;
      RECT 1.8550 1.3450 1.9800 1.5400 ;
      RECT 1.8800 0.5100 2.2400 0.6100 ;
      RECT 0.2650 1.6450 0.7450 1.7350 ;
      RECT 0.2650 1.2400 0.3550 1.6450 ;
      RECT 0.2350 0.9950 0.3550 1.2400 ;
      RECT 0.2650 0.7500 0.3550 0.9950 ;
      RECT 2.1000 1.4700 3.5750 1.5600 ;
      RECT 3.3300 1.4500 3.5750 1.4700 ;
      RECT 2.3800 0.4800 3.5650 0.5700 ;
      RECT 3.3900 0.4600 3.5650 0.4800 ;
      RECT 2.1000 0.8050 2.2000 1.4700 ;
      RECT 2.1000 0.7150 2.4700 0.8050 ;
      RECT 2.3800 0.5700 2.4700 0.7150 ;
      RECT 3.6850 1.3150 3.7850 1.5500 ;
      RECT 3.1900 1.2150 3.7850 1.3150 ;
      RECT 3.1900 1.0850 3.2900 1.2150 ;
      RECT 2.9050 0.9850 3.2900 1.0850 ;
      RECT 3.1900 0.7700 3.2900 0.9850 ;
      RECT 3.1900 0.6700 3.7900 0.7700 ;
      RECT 3.6800 0.4300 3.7900 0.6700 ;
      RECT 1.3050 1.4700 1.7450 1.5600 ;
      RECT 1.5900 0.8400 1.7950 0.9500 ;
      RECT 1.6550 1.5600 1.7450 1.6500 ;
      RECT 1.6550 0.9500 1.7450 1.4700 ;
      RECT 1.6550 1.6500 4.0150 1.7400 ;
      RECT 3.4600 0.8650 4.1350 0.9650 ;
      RECT 3.9150 1.1050 4.0150 1.6500 ;
      RECT 3.9150 0.8650 4.1350 1.1050 ;
      RECT 3.4450 1.9200 3.6550 1.9900 ;
      RECT 1.3950 1.9000 4.4300 1.9200 ;
      RECT 4.1650 1.9200 4.4300 1.9900 ;
      RECT 1.3950 1.8300 4.2700 1.9000 ;
      RECT 1.3950 1.7400 1.4850 1.8300 ;
      RECT 0.8550 1.6500 1.4850 1.7400 ;
      RECT 0.4550 0.9300 0.5450 1.4450 ;
      RECT 0.8550 1.5350 0.9450 1.6500 ;
      RECT 0.4550 1.4450 0.9450 1.5350 ;
      RECT 0.4550 0.8400 1.2800 0.9300 ;
      RECT 4.4150 1.3400 4.8600 1.4300 ;
      RECT 4.4150 0.7700 4.5150 1.3400 ;
      RECT 4.4150 0.6600 4.6250 0.7700 ;
      RECT 4.1400 1.5200 5.3850 1.6100 ;
      RECT 4.8150 0.6600 5.3700 0.7500 ;
      RECT 4.1400 1.6100 4.2600 1.6750 ;
      RECT 4.1400 1.2700 4.3250 1.5200 ;
      RECT 4.2250 0.7700 4.3250 1.2700 ;
      RECT 3.9150 0.6700 4.3250 0.7700 ;
      RECT 4.8150 0.7500 4.9050 1.0750 ;
      RECT 3.9150 0.4300 4.0750 0.6700 ;
      RECT 4.9700 1.1650 5.0600 1.5200 ;
      RECT 4.8150 1.0750 5.0600 1.1650 ;
      RECT 5.5650 1.0500 5.8550 1.1500 ;
      RECT 4.3900 1.7000 5.6550 1.7900 ;
      RECT 5.5650 1.1500 5.6550 1.7000 ;
      RECT 5.5650 0.5700 5.6550 1.0500 ;
      RECT 4.1700 0.4800 5.6550 0.5700 ;
      RECT 4.1700 0.4600 4.3950 0.4800 ;
  END
END ADDFH_X1P4M_A12TH

MACRO ADDFH_X2M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 6.2450 2.7200 ;
        RECT 2.6200 2.0450 2.7900 2.0800 ;
        RECT 3.1400 2.0450 3.3100 2.0800 ;
        RECT 4.9350 2.0350 5.1050 2.0800 ;
        RECT 5.4500 1.8700 5.6200 2.0800 ;
        RECT 6.0050 1.7600 6.1050 2.0800 ;
    END
  END VDD

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7700 1.2500 1.5650 1.3500 ;
        RECT 1.4650 1.0750 1.5650 1.2500 ;
    END
    ANTENNAGATEAREA 0.2451 ;
  END B

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 6.2450 0.3200 ;
        RECT 0.4000 0.3200 0.6100 0.3600 ;
        RECT 6.0050 0.3200 6.1050 0.6400 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6500 0.7600 2.7500 1.2500 ;
        RECT 2.6500 1.2500 3.0800 1.3800 ;
        RECT 2.6500 0.6600 3.0800 0.7600 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END CO

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7450 1.2500 6.1500 1.3500 ;
        RECT 5.7450 1.3500 5.8450 1.7150 ;
        RECT 6.0500 0.9500 6.1500 1.2500 ;
        RECT 5.7450 0.8500 6.1500 0.9500 ;
        RECT 5.7450 0.4300 5.8450 0.8500 ;
    END
    ANTENNADIFFAREA 0.325 ;
  END SUM

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6450 1.0500 1.1900 1.1600 ;
    END
    ANTENNAGATEAREA 0.0906 ;
  END A

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2350 0.9800 5.3900 1.2100 ;
        RECT 5.0100 0.8500 5.3900 0.9800 ;
    END
    ANTENNAGATEAREA 0.0975 ;
  END CI
  OBS
    LAYER M1 ;
      RECT 0.0450 0.4800 1.5550 0.5700 ;
      RECT 0.0450 1.4500 0.1750 1.8300 ;
      RECT 0.0450 0.8850 0.1350 1.4500 ;
      RECT 0.0450 0.5700 0.1750 0.8850 ;
      RECT 0.0450 1.8300 1.2750 1.9200 ;
      RECT 0.2650 0.6600 1.9800 0.7500 ;
      RECT 1.8900 0.7500 1.9800 1.3450 ;
      RECT 1.8800 0.6100 1.9800 0.6600 ;
      RECT 1.8550 1.3450 1.9800 1.5400 ;
      RECT 1.8800 0.5100 2.2400 0.6100 ;
      RECT 0.2650 1.6450 0.7350 1.7350 ;
      RECT 0.2650 1.2400 0.3550 1.6450 ;
      RECT 0.2350 0.9950 0.3550 1.2400 ;
      RECT 0.2650 0.7500 0.3550 0.9950 ;
      RECT 2.1000 1.4700 3.5750 1.5600 ;
      RECT 3.3300 1.4500 3.5750 1.4700 ;
      RECT 2.4000 0.4800 3.5650 0.5700 ;
      RECT 3.3400 0.4600 3.5650 0.4800 ;
      RECT 2.1000 0.8050 2.2000 1.4700 ;
      RECT 2.1000 0.7150 2.4900 0.8050 ;
      RECT 2.4000 0.5700 2.4900 0.7150 ;
      RECT 3.6850 1.3150 3.7850 1.5500 ;
      RECT 3.1900 1.2150 3.7850 1.3150 ;
      RECT 3.1900 1.0850 3.2900 1.2150 ;
      RECT 2.9050 0.9850 3.2900 1.0850 ;
      RECT 3.1900 0.7700 3.2900 0.9850 ;
      RECT 3.1900 0.6700 3.7900 0.7700 ;
      RECT 3.6800 0.4300 3.7900 0.6700 ;
      RECT 1.3050 1.4700 1.7450 1.5600 ;
      RECT 1.5900 0.8400 1.7950 0.9500 ;
      RECT 1.6550 1.5600 1.7450 1.6500 ;
      RECT 1.6550 0.9500 1.7450 1.4700 ;
      RECT 1.6550 1.6500 4.0150 1.7400 ;
      RECT 3.4250 0.8650 4.1350 0.9650 ;
      RECT 3.9150 1.1050 4.0150 1.6500 ;
      RECT 3.9150 0.8650 4.1350 1.1050 ;
      RECT 3.4400 1.9200 3.6550 1.9900 ;
      RECT 1.3950 1.9000 4.4400 1.9200 ;
      RECT 4.1550 1.9200 4.4400 1.9900 ;
      RECT 1.3950 1.8300 4.2600 1.9000 ;
      RECT 1.3950 1.7400 1.4850 1.8300 ;
      RECT 0.8550 1.6500 1.4850 1.7400 ;
      RECT 0.4550 0.9300 0.5450 1.4450 ;
      RECT 0.8550 1.5350 0.9450 1.6500 ;
      RECT 0.4550 1.4450 0.9450 1.5350 ;
      RECT 0.4550 0.8400 1.2800 0.9300 ;
      RECT 4.4150 1.3300 4.8600 1.4200 ;
      RECT 4.4150 0.7700 4.5150 1.3300 ;
      RECT 4.4150 0.6600 4.6300 0.7700 ;
      RECT 4.1400 1.5100 5.3900 1.6000 ;
      RECT 4.8150 0.6600 5.3900 0.7500 ;
      RECT 4.1400 1.6000 4.2600 1.6750 ;
      RECT 4.1400 1.2550 4.3250 1.5100 ;
      RECT 4.2250 0.7700 4.3250 1.2550 ;
      RECT 3.9150 0.6700 4.3250 0.7700 ;
      RECT 4.8150 0.7500 4.9050 1.0750 ;
      RECT 3.9150 0.4300 4.0750 0.6700 ;
      RECT 4.9700 1.1650 5.0600 1.5100 ;
      RECT 4.8150 1.0750 5.0600 1.1650 ;
      RECT 5.5650 1.0500 5.8550 1.1500 ;
      RECT 4.3700 1.6900 5.6550 1.7800 ;
      RECT 5.5650 1.1500 5.6550 1.6900 ;
      RECT 5.5650 0.5700 5.6550 1.0500 ;
      RECT 4.1700 0.4800 5.6550 0.5700 ;
      RECT 4.1700 0.4600 4.3950 0.4800 ;
  END
END ADDFH_X2M_A12TH

MACRO ADDF_X1M_A12TH
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 2.4 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.0450 -0.3200 4.2450 0.3200 ;
        RECT 0.3550 0.3200 0.4550 0.5800 ;
        RECT 1.8850 0.3200 1.9850 0.6300 ;
        RECT 3.7100 0.3200 3.8800 0.5050 ;
    END
  END VSS

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0900 1.6500 0.3900 1.7500 ;
        RECT 0.0900 0.4850 0.1900 1.6500 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END CO

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 0.9150 4.1500 1.2900 ;
        RECT 4.0150 1.2900 4.1500 1.7100 ;
        RECT 4.0150 0.4950 4.1500 0.9150 ;
    END
    ANTENNADIFFAREA 0.284375 ;
  END S

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8300 0.8500 3.6800 0.9500 ;
        RECT 0.8300 0.9500 1.0400 1.0100 ;
        RECT 3.5800 0.9500 3.6800 1.2800 ;
    END
    ANTENNAGATEAREA 0.3138 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0450 2.0800 4.2450 2.7200 ;
        RECT 3.7100 1.8950 3.8800 2.0800 ;
        RECT 2.4050 1.8550 2.5050 2.0800 ;
        RECT 0.3500 1.8400 0.4500 2.0800 ;
        RECT 0.8850 1.7700 0.9850 2.0800 ;
        RECT 1.8850 1.7700 1.9850 2.0800 ;
    END
  END VDD

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9350 1.2500 3.2600 1.3500 ;
    END
    ANTENNAGATEAREA 0.2217 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4650 1.1000 3.4700 1.1500 ;
        RECT 1.1800 1.0500 3.4700 1.1000 ;
        RECT 0.4650 1.1500 1.2800 1.2000 ;
    END
    ANTENNAGATEAREA 0.3138 ;
  END A
  OBS
    LAYER M1 ;
      RECT 0.6300 1.5900 1.2050 1.6800 ;
      RECT 1.1150 1.6800 1.2050 1.8300 ;
      RECT 1.1150 1.8300 1.7400 1.9200 ;
      RECT 1.5700 1.6300 1.7400 1.8300 ;
      RECT 0.6300 1.6800 0.7200 1.9800 ;
      RECT 0.5700 0.4800 1.7600 0.5700 ;
      RECT 2.1450 1.6200 2.7950 1.7100 ;
      RECT 2.6950 1.7100 2.7950 1.9900 ;
      RECT 2.1450 1.7100 2.2450 1.9900 ;
      RECT 2.0900 0.4800 2.8600 0.5700 ;
      RECT 1.3100 1.4700 2.9550 1.5300 ;
      RECT 0.2800 1.4400 2.9550 1.4700 ;
      RECT 1.3100 1.5300 1.4800 1.6850 ;
      RECT 0.2800 1.3800 1.4800 1.4400 ;
      RECT 0.2800 0.6700 1.5000 0.7600 ;
      RECT 0.2800 0.7600 0.3700 1.3800 ;
      RECT 2.9550 1.7000 3.9050 1.7900 ;
      RECT 3.8150 0.6850 3.9050 1.7000 ;
      RECT 2.9950 0.5950 3.9050 0.6850 ;
      RECT 2.9550 1.7900 3.1250 1.9900 ;
      RECT 2.9950 0.4400 3.0950 0.5950 ;
  END
END ADDF_X1M_A12TH
  
END LIBRARY
